// Matrix that loads data from the given memory / hardcoded for our multiplications

module matrix(input logic[9:0] counter1, input logic[6:0] counter2,
			output shortint counter1_out[0:99], counter2_out[0:9],
			output shortint counter1_bias[0:99], counter2_bias[0:9]);
			
	assign counter1_bias = '{0,0,0,1,0,-2,1,-1,-1,-2,0,0,0,-1,3,-1,2,0,1,3,-2,1,-3,2,-2,0,2,2,1,-3,1,-1,1,1,-1,-2,-2,-1,0,0,-1,-2,1,-1,0,0,-3,-1,-3,-4,-1,-1,1,2,-1,0,3,-1,1,0,-1,1,-1,-1,0,-1,0,0,-1,-4,0,0,-3,-3,-2,2,-1,0,-1,-2,-2,3,0,0,-2,-2,-1,-4,0,-1,-2,-1,-1,-1,0,1,-3,0,-3,1};
	assign counter2_bias = '{-3,-2,0,-2,-3,-2,-2,-3,-1,-2};
	
			
	always_comb
	// Combination Block for counter1 matrix
	begin
		case (counter1)
			default: counter1_out = '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
			0: counter1_out = '{0,1,1,0,-2,-1,0,2,0,0,0,-1,-1,0,0,1,0,0,0,0,0,0,0,0,1,1,1,-1,0,-1,1,0,1,-2,-1,-2,0,0,-2,0,1,-1,0,0,1,-1,0,0,0,1,1,-1,-1,0,1,1,1,1,0,0,0,-2,0,0,-2,-1,-2,-1,-1,-1,-1,0,1,-1,0,1,-2,2,0,0,1,1,0,1,0,-2,1,0,0,1,1,2,-1,-1,0,-1,1,-1,-1,0};
			1: counter1_out = '{1,0,-1,2,0,1,1,-1,0,1,1,1,0,-1,0,-1,-1,-1,-1,1,-1,1,1,0,0,-1,0,0,-1,-3,1,0,-2,0,0,0,1,1,-3,0,1,0,-1,0,-1,1,0,0,-3,2,0,-1,1,0,0,-1,0,-1,2,0,-2,2,1,1,-1,0,-1,0,2,-1,1,-3,0,-1,0,1,2,1,-1,0,3,0,1,-3,0,-2,0,0,0,1,-1,0,0,0,0,0,-1,2,-1,1};
			2: counter1_out = '{-2,-1,0,-1,0,-1,-2,0,-2,-3,-1,1,0,-1,0,1,1,0,2,0,-1,0,-1,-2,0,0,0,-1,-2,0,-1,0,-1,-1,0,0,-2,-1,1,-1,-1,2,1,1,0,-1,1,-1,-2,0,1,-2,-1,-1,-1,1,-1,-1,0,1,-1,1,0,0,0,0,-1,0,1,0,0,1,0,2,-3,-1,0,-1,0,-1,1,-2,-1,-1,-1,0,0,-1,0,-1,-3,-2,1,1,0,1,-1,1,1,1};
			3: counter1_out = '{-1,-2,1,-2,-1,1,0,1,0,-1,0,1,1,-1,-2,0,0,0,1,0,0,-2,1,0,0,-1,1,-1,-1,0,1,0,0,0,2,-1,0,1,1,-1,0,1,0,2,-1,-1,-1,0,2,-1,1,-1,-1,-1,-1,-2,1,-1,2,1,0,1,1,2,0,0,0,0,0,-1,0,-1,0,0,0,-1,-2,1,1,1,1,1,-1,-1,1,1,-1,0,1,0,0,2,-1,0,0,0,-2,0,1,-1};
			4: counter1_out = '{3,-2,0,0,1,2,-1,0,-1,1,0,-2,0,-1,-1,1,1,0,2,-1,-1,-1,0,-1,-2,-1,0,1,0,-1,1,2,1,0,0,-1,0,1,2,1,-2,1,1,-1,-1,0,0,2,1,1,-1,0,2,-1,0,-1,1,0,1,-1,-2,0,0,1,-1,0,-2,0,1,0,0,0,1,-1,-3,-2,0,-1,-1,1,1,0,0,1,-2,2,2,1,-1,2,2,0,3,0,0,0,-1,-1,0,0};
			5: counter1_out = '{-1,0,0,0,0,1,-1,0,1,0,-1,0,0,1,0,1,3,1,0,-1,0,-1,-1,-1,0,1,0,0,0,0,0,-1,0,0,0,0,-1,0,2,1,1,1,1,-1,-1,1,1,1,1,0,2,1,-3,0,0,1,-1,-1,-1,0,0,1,-1,0,0,1,2,-1,-1,0,0,2,0,-1,0,-2,0,-2,0,-1,1,-1,1,0,1,0,1,0,-1,-1,1,-1,0,-1,-1,2,0,-1,1,1};
			6: counter1_out = '{2,1,1,1,1,0,2,0,0,0,0,-1,0,1,0,-1,0,1,-1,1,0,-2,-2,1,-3,0,1,1,-1,-1,1,-1,0,1,-1,0,0,0,-1,0,1,0,1,2,0,1,0,0,-2,-1,0,1,0,-1,0,1,1,0,0,1,-1,0,0,1,-3,-1,0,0,-1,0,-1,0,0,-1,0,0,1,0,0,-1,-1,-1,0,1,0,1,-1,-1,2,0,1,1,0,1,0,0,-1,0,-1,-1};
			7: counter1_out = '{0,-1,1,0,0,1,2,0,1,1,-2,0,1,-1,2,1,-1,1,1,-1,1,2,-1,0,-1,1,-1,-1,2,0,2,1,1,-1,2,-1,-1,-1,0,0,-2,0,-1,2,0,-1,1,0,0,-2,0,0,1,0,1,0,2,1,0,0,1,2,1,-2,-1,-1,1,1,0,0,-1,-1,2,2,1,1,0,0,0,-1,0,-3,0,0,2,1,0,0,-1,0,-2,-1,-1,1,-1,-1,0,1,-1,0};
			8: counter1_out = '{0,0,0,-1,0,-1,0,0,1,1,-1,0,1,0,0,0,-1,-1,-1,1,0,0,1,-1,0,0,0,-1,0,-1,0,0,1,0,1,-2,-2,1,1,0,-1,0,1,-1,-1,2,1,0,0,0,-1,0,0,1,1,1,-1,0,0,0,1,1,0,0,2,0,0,0,-1,1,-1,-2,0,0,0,-2,0,-1,0,0,0,0,0,0,1,0,0,0,1,1,2,-1,-1,0,1,-1,-1,-1,-1,-2};
			9: counter1_out = '{1,1,-1,1,0,-1,0,0,2,0,-1,0,-1,2,2,-2,-1,0,0,0,0,1,-1,-2,0,0,0,0,0,2,1,-1,0,0,0,-1,0,-1,-1,-2,-1,0,0,-1,1,-1,2,1,-1,-2,1,1,1,1,2,-2,1,0,0,-1,0,2,0,0,1,1,1,-1,0,0,0,0,1,2,1,0,-1,0,0,1,0,-1,-1,-1,-1,0,0,1,0,-1,0,0,-1,0,0,0,0,-1,1,0};
			10: counter1_out = '{0,1,-1,1,-1,-1,0,1,0,1,-2,0,-1,1,0,-3,1,2,2,0,-1,2,0,1,-1,0,-1,1,1,0,1,0,-2,0,1,-1,1,1,-1,0,1,0,-1,0,0,-2,0,1,0,0,-1,-1,0,-1,2,1,1,1,-1,-1,-1,1,-1,-1,0,-1,-1,0,0,0,-1,0,-2,-2,1,-1,0,1,1,0,1,0,1,0,-1,-1,1,-1,0,0,1,1,0,0,0,0,0,0,0,0};
			11: counter1_out = '{0,0,0,-1,-1,1,2,-1,0,-1,0,0,0,0,0,1,0,1,0,1,0,-1,0,1,0,0,0,0,0,0,1,1,-1,2,1,-1,1,0,-1,0,0,-1,-1,-1,1,1,0,0,0,-2,1,1,-1,1,0,-1,0,1,0,-1,-1,-1,1,-1,-1,0,0,-1,0,-1,0,-1,-1,0,1,0,-1,-1,-1,-1,-1,0,-2,-1,-1,-2,0,-1,1,-1,0,-1,0,0,0,0,0,0,0,0};
			12: counter1_out = '{-1,-1,1,-2,0,0,1,0,-1,1,-2,-2,1,1,-1,-2,-2,-1,-1,-1,-1,-1,0,-1,1,0,-1,-2,0,1,-1,0,0,-1,0,0,0,-2,2,0,0,1,0,0,1,-1,0,0,0,-1,1,0,-2,-1,-1,0,0,-1,0,0,-1,0,0,0,0,0,2,0,-2,0,0,0,0,0,-2,-1,1,0,1,-1,0,0,0,0,-1,-1,0,0,0,0,-1,1,1,0,0,-1,2,0,0,-1};
			13: counter1_out = '{-1,1,-1,-1,0,0,-1,0,0,0,-1,0,-2,1,0,0,1,1,-1,0,1,0,0,1,-1,1,1,2,0,1,-1,-2,1,-1,2,0,-1,-1,1,-1,1,-1,-1,-2,0,1,1,1,-1,0,0,0,0,0,-1,0,0,1,0,0,-1,0,1,0,-2,0,0,0,0,1,0,-1,-2,-1,2,-1,-1,0,2,1,1,1,-2,0,-1,1,1,-2,-1,0,1,1,0,-1,0,1,1,-2,0,-1};
			14: counter1_out = '{2,-1,-1,-1,-1,0,0,0,1,-2,0,0,-2,1,0,1,1,-1,2,2,1,0,0,-1,0,-1,1,-1,-1,1,2,2,-1,1,-1,-1,-1,0,0,0,-1,2,-1,0,-1,-2,1,2,1,1,0,-1,0,0,0,1,1,2,2,0,-1,-1,2,0,1,0,0,2,0,-1,0,0,1,1,2,-3,1,0,-2,-2,0,0,0,2,-3,-1,1,0,1,1,-1,0,-1,0,1,0,0,0,1,-1};
			15: counter1_out = '{0,0,0,1,-1,0,0,1,2,-1,0,-1,1,0,1,1,0,0,1,-2,0,-1,0,1,-1,-1,1,1,0,0,-1,-1,1,0,0,0,0,-1,-1,1,0,0,-1,-2,0,-1,-2,1,1,0,1,0,1,0,-1,0,-1,1,0,-2,1,1,0,-1,0,0,1,1,1,1,1,1,0,-1,0,1,2,1,1,0,-1,1,2,-1,-1,0,1,-1,-1,-1,0,0,1,-1,1,1,-1,0,1,0};
			16: counter1_out = '{0,-1,0,0,0,3,-1,0,0,-1,1,-1,0,1,-1,0,-1,0,0,0,-2,0,0,0,-1,-1,-1,0,-1,-1,0,0,0,1,-1,0,-1,1,0,0,0,1,0,1,-1,-2,2,0,1,0,-1,-2,-1,0,0,-1,1,1,0,-1,-1,0,1,1,-1,0,0,1,0,0,0,0,1,-1,1,-1,2,0,2,0,2,0,2,-1,-1,-1,-1,0,-1,-1,2,1,1,0,1,0,0,1,1,2};
			17: counter1_out = '{0,0,1,-1,1,-1,0,-1,0,-2,-1,0,0,2,0,-1,-2,-1,-1,-2,0,1,-1,0,-1,0,0,-1,-1,1,1,0,-1,2,1,0,0,1,-1,-1,0,1,2,0,-1,0,1,2,-2,0,0,0,0,-1,0,0,-2,0,0,1,0,1,1,0,0,0,2,0,-1,-1,-1,3,1,1,1,-1,0,0,0,0,1,1,-1,0,1,1,0,-1,2,0,1,1,1,1,-1,1,2,0,1,0};
			18: counter1_out = '{-1,-1,-2,0,0,1,1,1,0,2,0,2,-1,-2,0,-1,1,1,-1,-1,0,2,1,-1,0,-1,2,0,0,1,0,0,0,0,3,1,0,-1,0,-1,-1,1,0,-1,-2,1,-1,0,1,3,-2,-1,1,0,-1,1,-1,2,0,0,0,1,-1,-1,-2,1,-1,0,0,1,-1,0,1,3,-2,2,-1,1,0,2,1,-2,1,-1,2,0,-1,2,0,1,1,0,0,1,2,0,0,2,-2,1};
			19: counter1_out = '{0,2,-1,0,-2,0,-1,-2,1,-2,-1,1,0,-1,0,-1,1,0,-3,1,-1,-1,0,1,-2,-1,0,-1,0,1,-1,-2,-2,0,1,1,1,0,0,1,0,2,1,-2,0,1,-1,0,0,1,-1,1,-1,0,-2,-2,1,-1,0,1,-2,1,0,1,0,-1,0,0,-2,0,1,0,-2,0,1,0,-1,1,2,1,0,0,0,-1,-1,0,0,0,-1,-1,2,-1,0,-1,0,-2,1,0,2,1};
			20: counter1_out = '{1,-1,-1,1,-1,1,0,-1,1,0,1,0,0,1,1,1,-2,0,-2,2,1,0,0,0,-1,2,0,0,0,-1,2,-2,1,0,-1,1,0,0,0,0,1,-1,0,0,-1,-1,0,-2,0,1,-1,1,-2,0,0,-1,-1,0,0,0,1,-1,1,2,0,1,0,-1,0,1,0,1,1,0,0,2,-1,-3,0,-1,-1,1,0,0,0,1,0,0,1,1,-1,2,0,0,0,1,-1,1,1,-1};
			21: counter1_out = '{0,-1,0,1,0,-1,1,-1,1,2,-3,1,0,0,1,2,0,-1,-2,-1,-1,-1,1,-1,-2,0,0,-1,-1,1,0,-2,0,0,0,0,0,0,0,0,1,-1,-1,0,1,0,-1,0,-2,0,1,0,-1,-1,1,-1,-1,0,-2,-2,0,0,0,0,0,-2,-1,0,-1,0,0,0,1,0,2,2,-2,-1,1,1,-1,1,0,-1,2,0,0,0,-1,-2,-1,1,-1,2,0,0,-2,0,-1,2};
			22: counter1_out = '{0,-2,1,0,1,1,-1,2,0,0,0,1,0,0,0,0,-2,-1,-1,1,1,-1,0,1,-1,-1,0,0,0,-2,-1,-2,-1,0,-1,0,0,0,1,2,1,-2,0,1,0,1,1,2,0,0,1,0,1,0,-2,-1,2,-1,-1,2,0,0,-2,-1,0,-2,1,-1,-2,0,0,-1,-2,0,1,-1,-2,-1,0,1,-1,-1,1,-1,-1,1,0,0,0,2,2,-1,1,0,1,-1,0,1,0,-1};
			23: counter1_out = '{2,-1,1,-1,-1,-1,0,2,2,0,1,-1,1,1,0,-1,-1,0,0,-1,0,-1,-1,-1,1,1,0,-1,0,1,-3,0,-1,2,-2,0,-1,0,0,-1,1,1,-1,1,-1,0,1,0,0,0,-1,0,0,-1,2,0,0,-3,-2,0,0,2,2,-1,-1,1,0,1,-1,1,1,1,-1,-1,0,0,1,0,1,2,2,0,0,1,2,0,0,-1,0,1,2,2,0,2,1,-1,1,0,0,0};
			24: counter1_out = '{0,0,0,0,2,0,0,0,-1,0,0,0,0,0,0,-1,0,-1,-1,0,0,2,0,0,-1,-1,-1,-1,1,0,2,0,1,1,0,-2,-1,0,-2,1,-1,-1,-1,-1,0,0,0,1,0,1,0,0,1,0,2,0,2,0,0,0,0,1,-1,-1,1,0,2,0,0,0,0,1,-1,-1,1,-1,-1,0,0,1,-1,-1,0,0,1,-1,1,0,0,0,-1,-1,0,1,1,0,-1,0,1,0};
			25: counter1_out = '{1,0,1,0,1,1,2,0,1,0,0,-1,0,0,-1,0,0,0,0,-2,0,1,-1,1,-1,1,0,0,-1,0,-1,1,1,0,0,-1,0,1,0,1,-1,0,-1,-2,0,-2,0,1,0,1,1,2,0,1,0,1,-2,-2,0,0,0,0,-1,2,2,0,2,0,1,-1,0,1,1,0,0,0,0,-1,-1,-1,2,1,1,-2,-1,1,2,0,1,1,0,1,1,1,1,0,-1,1,-1,0};
			26: counter1_out = '{0,0,0,1,-1,-2,1,-1,1,2,0,0,0,0,-2,0,2,1,-2,-1,0,1,1,2,1,0,0,1,0,0,1,1,-1,-1,0,0,-1,0,2,-3,0,1,0,-1,0,1,1,1,2,-1,0,1,-1,1,1,1,1,-1,0,-1,1,1,1,-1,1,-1,0,0,0,0,0,0,0,-1,-1,-1,0,-1,1,0,1,0,-1,-2,-2,0,1,1,-1,-1,-2,0,1,1,1,-1,1,0,0,0};
			27: counter1_out = '{0,0,-2,1,0,-1,0,0,1,1,0,1,-1,0,0,1,0,0,0,-1,1,1,1,1,-1,-2,-1,-1,0,1,-1,1,0,1,0,-1,-1,1,-1,1,0,2,0,0,2,0,1,0,0,1,0,-1,-1,-1,1,0,0,-1,-1,2,0,0,1,1,-1,-1,1,0,0,-1,-1,-1,-1,1,1,1,0,0,0,1,2,1,1,0,-1,-2,0,-1,2,1,2,1,0,0,1,0,0,-1,0,1};
			28: counter1_out = '{1,0,0,0,1,1,0,0,-1,0,0,-1,-1,0,0,-1,-3,-1,-1,1,1,0,1,-2,0,-2,1,0,-2,1,0,2,-1,1,-2,1,1,0,1,2,-1,-1,-1,0,1,1,-1,0,0,0,1,0,0,1,0,-1,0,-2,-1,-3,1,1,1,-1,1,0,1,1,-1,1,-1,-2,0,1,1,-1,0,2,1,-3,0,2,1,1,0,1,-1,0,0,-1,0,-1,-1,1,-2,-1,0,1,1,0};
			29: counter1_out = '{-1,0,2,1,-1,-2,-2,-2,-2,0,-2,0,0,0,1,-2,1,-1,-2,-1,0,0,-1,0,2,0,1,1,1,-1,0,2,1,2,2,-1,0,0,1,0,1,2,-1,0,0,0,0,-1,0,0,0,0,2,0,-2,2,-1,0,-1,1,0,1,0,1,-1,0,0,0,0,-1,0,0,1,1,-1,1,-1,0,2,-2,0,-1,1,1,2,0,2,0,-1,2,1,1,0,0,-1,0,0,1,0,0};
			30: counter1_out = '{-1,1,1,1,-1,-1,0,-2,-2,0,0,1,-1,1,0,-3,0,1,0,1,-2,2,-2,1,0,-2,1,2,0,-1,-1,0,0,0,0,1,-2,-2,0,0,0,-1,-1,0,0,-1,1,1,1,0,0,0,0,1,0,-1,-2,-1,0,2,-1,1,-1,0,0,0,-1,0,0,0,-1,2,2,-1,-2,0,-1,2,-1,1,0,1,0,1,-1,0,-2,0,-1,1,1,-1,0,0,-1,2,0,-2,-1,-2};
			31: counter1_out = '{-1,0,1,0,1,0,0,1,0,-1,0,1,0,-1,2,1,2,-1,0,0,-1,1,-1,1,0,0,1,1,0,1,0,-2,-1,-1,-1,-1,0,-1,0,1,0,1,-1,0,1,-1,-1,1,-1,1,0,0,1,-1,1,0,2,1,0,2,-1,0,-1,0,-2,2,-1,0,1,2,0,1,0,1,0,0,1,0,-1,0,-2,1,0,0,-1,1,0,1,0,1,1,0,1,-1,0,1,0,-1,1,-1};
			32: counter1_out = '{1,-1,1,0,-1,0,1,1,1,2,1,-1,-1,3,0,-1,1,-1,-1,-1,0,0,1,0,0,0,0,0,2,-1,-1,-1,-1,1,1,1,2,0,-1,1,0,1,1,-1,-1,0,-1,0,1,0,0,-1,0,0,0,-1,1,-1,-2,0,-3,1,-1,0,0,-2,1,-1,0,-1,1,1,0,1,0,-1,-1,0,0,0,1,2,0,0,-2,1,0,-2,-1,-1,2,-1,-1,0,-1,0,1,-1,0,0};
			33: counter1_out = '{-1,-1,1,1,0,2,1,-1,-1,1,0,-1,0,0,1,0,1,1,0,1,2,0,0,-2,-2,0,1,2,-1,-2,0,0,-2,1,-1,-1,-2,0,-1,0,-1,-1,1,0,1,2,0,0,1,1,1,0,0,-1,2,2,1,-1,-1,-1,1,1,0,1,-1,1,1,-2,1,-2,-2,0,-1,-1,0,1,0,1,-1,0,0,0,2,2,0,-1,-2,-2,0,-1,0,-1,1,1,-1,-1,-1,0,0,1};
			34: counter1_out = '{-1,1,-1,1,0,-2,-1,2,1,0,0,0,-1,1,0,0,0,0,0,-2,0,0,2,2,1,0,0,0,1,-1,1,1,0,-2,1,0,-1,0,1,-1,-1,-1,-1,-1,0,0,0,2,0,0,2,-2,0,0,-1,-1,0,1,-1,1,-2,0,0,-1,-1,0,1,-1,1,1,0,0,0,0,0,0,1,2,-1,1,1,1,-1,-1,0,-1,-1,-3,0,0,-1,-1,-1,0,-1,0,0,0,-2,1};
			35: counter1_out = '{-1,0,-1,-1,0,1,0,-1,1,0,1,-2,0,0,0,-1,0,-2,1,2,0,-1,-2,2,1,1,0,0,0,0,-1,2,-1,0,1,0,-1,1,1,2,-2,-1,-2,-1,4,0,0,-1,1,2,0,1,0,1,-1,-1,2,1,0,1,-1,-1,0,-1,0,1,0,0,0,-1,-1,0,0,-1,0,-2,-1,0,0,-2,0,-1,1,-1,-1,0,0,-1,0,0,2,0,0,-2,1,2,0,3,-1,0};
			36: counter1_out = '{1,-1,-1,-1,1,0,1,0,-1,0,-2,0,-1,0,-1,3,1,0,1,1,-1,-1,2,-1,0,1,1,-1,0,0,1,0,2,-1,0,0,0,0,-1,0,-1,0,0,2,2,0,1,-2,1,0,1,0,-1,0,1,0,-1,-1,-1,1,-2,-1,0,0,0,2,0,0,1,0,0,-1,-1,0,0,1,0,0,1,0,1,-1,-1,-1,-1,0,0,0,-1,0,-1,1,0,0,0,0,2,1,1,0};
			37: counter1_out = '{-1,1,0,1,1,1,1,1,1,0,0,0,1,0,2,1,1,1,-1,-1,-1,1,1,0,0,0,0,0,-2,-1,1,1,-2,2,0,0,0,-1,1,-1,1,-1,1,0,0,0,-1,-1,0,-1,1,0,1,0,1,1,-1,0,-1,0,-1,1,1,-1,0,0,1,0,0,-1,0,0,0,0,0,0,-2,0,-1,-1,0,3,-1,-1,-1,0,-1,0,1,0,0,-1,-1,1,1,0,0,2,-1,-2};
			38: counter1_out = '{2,0,0,-2,1,1,0,-1,-1,-2,0,1,0,0,1,0,1,2,2,-1,1,0,0,0,1,-2,-1,0,0,-1,-1,-2,0,0,-2,-1,1,1,-1,1,0,0,-1,0,0,-2,-1,0,0,-1,0,0,-1,0,-2,0,-1,-1,-2,1,-1,0,-1,1,0,-1,1,-1,-1,0,1,1,0,1,0,0,-1,-1,1,1,1,0,-1,0,0,0,1,-1,0,-1,-1,0,1,1,-1,0,-1,0,0,0};
			39: counter1_out = '{-2,-1,-1,-1,-1,1,-1,0,0,0,0,-1,0,0,-2,-1,0,0,0,-1,0,0,0,-2,1,0,-1,0,1,1,1,-1,-1,1,-1,0,0,0,1,0,1,0,0,1,0,-1,-1,-1,0,0,-1,0,-3,1,0,-1,-1,1,0,0,-1,1,-1,0,-2,0,-1,1,0,0,0,1,1,1,-1,0,0,0,0,0,0,0,1,1,0,2,1,-1,0,-1,0,0,0,0,0,1,0,-1,0,-1};
			40: counter1_out = '{-1,-1,-1,1,1,1,0,1,1,0,-1,-1,0,0,0,0,0,-1,-2,0,-2,4,0,-3,1,2,-1,2,0,2,2,0,-1,-1,0,1,1,0,2,-1,0,2,2,2,-1,1,0,-1,1,0,0,-1,-1,0,1,-2,1,1,-1,0,0,-2,-1,1,-1,-1,-2,0,-1,-1,1,0,1,0,-1,1,-1,2,0,0,0,-1,2,0,0,0,1,0,-1,0,1,-1,0,-1,0,-1,2,-2,1,-1};
			41: counter1_out = '{1,1,0,0,-2,-2,1,2,0,0,-2,2,0,0,2,0,1,0,0,-2,0,-1,-1,0,2,0,-2,0,-1,0,0,-1,-1,-2,1,0,0,1,0,1,1,-1,0,0,2,0,-1,0,0,-2,-1,1,0,0,-1,1,-2,0,-1,-1,0,2,-1,-1,-1,0,1,-1,0,-1,0,1,3,-1,0,0,0,1,0,0,0,-1,0,0,0,1,0,-1,0,1,1,1,1,0,1,0,-2,0,-1,1};
			42: counter1_out = '{0,0,0,-1,1,0,-1,-1,1,-1,1,2,1,0,1,-1,1,0,-1,0,1,-1,1,0,0,-1,0,0,-1,0,1,-2,-1,0,2,1,0,0,-1,1,1,0,-1,-2,-1,1,0,1,-1,1,-2,1,0,-1,-1,1,1,0,1,0,0,0,0,0,-1,0,1,0,0,0,1,1,-1,-1,-1,2,0,0,1,-1,1,1,-1,0,1,0,1,1,-2,1,1,2,-1,1,1,1,1,0,-1,-1};
			43: counter1_out = '{0,0,0,-1,2,-2,0,0,-1,0,-1,-2,1,-1,0,1,1,1,0,0,-1,-2,1,-1,-1,1,-1,0,0,0,0,0,-1,-1,0,-1,-2,-1,0,1,0,-1,0,0,0,-2,-1,2,0,2,2,-2,1,1,-1,-1,-1,-1,-1,0,0,0,0,1,0,-1,1,0,0,0,2,0,1,1,1,1,-2,1,0,2,-1,1,-1,0,2,0,1,0,-2,0,0,0,1,0,0,0,1,-1,0,2};
			44: counter1_out = '{1,-1,1,-1,0,-2,1,1,2,0,-1,1,1,1,-1,0,1,0,-1,0,-1,-1,0,1,-2,2,-1,0,-1,0,1,-1,-2,0,1,-3,0,-1,0,0,1,0,-1,-1,-1,1,-2,1,-1,1,0,-1,1,0,2,0,1,0,1,0,0,0,1,2,-1,1,2,-1,-2,1,1,-1,0,2,0,1,0,-1,0,0,1,-1,-1,1,0,-2,0,-1,2,-2,0,0,-1,0,0,-1,0,0,-1,-1};
			45: counter1_out = '{-1,0,0,-1,0,1,0,0,0,0,0,1,1,-1,-2,0,0,-1,0,0,0,1,0,-1,0,0,1,-1,0,0,1,-1,0,0,0,2,-1,2,-2,0,-1,0,-1,-1,0,0,0,0,2,-1,1,0,0,1,1,0,-1,0,0,0,0,0,-2,1,0,0,0,1,1,1,1,0,0,-1,2,0,0,-1,-1,-2,-1,0,-1,-1,0,0,0,-1,0,0,1,0,2,0,2,1,1,1,2,1};
			46: counter1_out = '{-1,-1,-1,-1,1,1,-1,1,-1,0,0,0,-1,1,0,0,1,0,-1,0,1,-2,0,0,2,-2,0,2,0,0,1,1,1,1,0,2,2,1,0,0,-1,0,0,-1,-2,2,0,-1,0,-1,0,2,0,0,0,0,-1,1,0,0,0,1,-1,1,0,0,2,-1,0,0,-2,1,0,0,0,0,-1,0,0,-2,0,0,-2,0,0,1,2,2,1,1,0,-1,0,-1,1,0,0,2,0,-1};
			47: counter1_out = '{0,-1,-1,-1,0,0,0,2,-1,0,-2,-1,0,-1,-1,-1,1,0,0,-1,0,1,0,1,-1,-1,-2,0,0,1,1,1,-2,0,0,1,-1,2,0,-2,0,0,0,0,0,1,-1,-1,-2,-1,2,-1,1,0,-1,-2,-1,0,-1,0,-2,0,0,-1,0,0,0,0,2,-1,-2,-1,0,1,2,-1,1,-1,1,-1,1,1,1,0,-1,-1,-1,0,-1,-1,0,-1,-1,1,0,-1,1,-1,0,1};
			48: counter1_out = '{-1,1,0,1,0,1,-1,-1,1,-1,-1,-1,-1,0,0,0,1,0,1,-1,1,0,1,1,-2,0,1,0,1,1,0,-1,1,0,0,0,-1,1,-1,1,0,1,-2,0,0,-2,0,-1,2,-1,0,0,0,0,-1,-1,-1,1,1,0,-1,0,0,-1,-1,-1,2,-2,0,0,2,-1,0,0,-2,0,1,-2,-1,-1,-1,0,-1,3,0,0,1,0,2,0,-1,-1,0,-1,1,-1,-1,0,0,0};
			49: counter1_out = '{-1,-1,-1,1,0,1,0,-1,-1,1,0,-2,0,1,0,2,0,0,0,0,-1,0,-2,-1,-1,2,0,-1,1,-1,0,0,0,-1,0,1,0,0,0,0,0,0,1,3,1,0,0,-2,0,1,0,-1,-1,-1,1,-1,0,2,0,0,1,0,0,-1,0,0,-1,0,-2,-1,0,1,1,1,1,-1,-1,-2,0,0,-2,-1,1,1,0,-1,-3,-1,-1,2,0,0,1,1,0,1,-1,0,-1,-1};
			50: counter1_out = '{-3,-1,0,0,0,-1,-1,0,1,1,1,2,-1,-1,1,-1,-1,1,-2,-2,0,-1,0,0,0,0,2,1,-2,-2,1,1,-1,0,0,0,2,0,-1,2,1,0,0,1,-1,-1,-2,0,-1,0,2,1,2,0,-1,0,0,-1,1,1,2,-1,-2,0,-1,0,1,0,-1,-1,-1,1,0,0,1,0,0,3,0,-2,2,-1,1,1,2,2,-1,0,-1,0,0,0,-1,0,-1,1,-1,-1,0,2};
			51: counter1_out = '{0,0,2,0,0,0,0,-2,1,1,-1,1,0,-1,0,-1,0,0,-1,-1,0,-1,0,0,0,0,-1,1,1,-1,-2,1,-1,1,0,1,1,1,0,3,0,0,-1,-2,0,0,-2,0,1,0,0,-1,0,-2,0,0,0,1,-1,0,1,-1,-2,2,1,0,0,0,1,0,0,0,-1,-1,0,0,-1,-1,1,0,1,-1,-2,1,0,1,0,-1,-1,1,0,1,-2,1,2,-1,-1,1,0,-2};
			52: counter1_out = '{1,0,0,1,1,1,0,-1,-1,-1,0,2,0,0,2,-1,1,1,0,0,-1,-1,0,0,-1,1,-1,0,-1,0,0,-1,1,-2,3,0,-1,-1,1,0,1,-1,0,0,1,2,0,1,0,2,-1,1,1,0,-1,0,1,0,0,0,1,-1,2,1,-1,-2,-2,1,-1,0,0,2,0,1,0,0,-1,1,0,2,0,3,-1,-1,0,0,-1,1,0,-1,0,-1,0,1,0,1,2,-1,0,0};
			53: counter1_out = '{1,2,0,0,1,1,0,1,0,0,1,-1,-1,0,0,0,1,-1,1,1,-1,0,-1,-2,1,3,0,-2,-1,0,-1,-1,-1,3,1,0,-1,0,0,0,1,-1,1,0,0,0,1,2,0,0,1,0,0,1,0,-1,2,0,0,1,1,0,0,1,1,0,-1,-1,2,1,-1,2,0,1,0,0,-1,-1,-1,0,0,0,2,0,1,0,0,1,-2,0,-1,-1,-1,-1,0,-2,0,-1,-2,-2};
			54: counter1_out = '{-1,0,-1,-2,1,0,-1,-1,0,-1,0,0,0,0,-1,-1,0,0,1,-1,-1,-1,1,-1,0,0,1,1,-1,0,2,0,0,0,0,0,0,-2,0,0,1,1,0,0,-1,3,0,1,1,0,0,-1,-1,0,2,1,0,1,-1,-1,-2,0,-1,1,0,1,1,0,0,1,0,1,-2,-2,1,1,1,0,-1,0,1,0,2,-1,1,-1,-1,1,0,-1,-1,0,-1,-1,1,1,-1,-1,-1,-1};
			55: counter1_out = '{0,1,0,1,0,-1,-1,0,1,-1,-1,0,1,1,0,0,0,1,0,2,-1,0,1,-1,0,-2,1,-2,-1,-1,-1,-1,0,1,0,0,1,0,0,0,0,1,0,0,-1,1,-1,1,2,2,0,-2,0,0,-1,0,0,1,0,-1,2,0,1,2,0,0,1,2,1,1,-1,1,1,1,0,0,1,-1,-1,2,1,0,0,0,0,1,1,-1,-1,-1,-1,-2,2,0,0,-1,0,1,1,-1};
			56: counter1_out = '{0,-2,-2,0,0,0,0,0,-1,-1,-1,0,2,2,1,1,2,0,-2,-1,0,1,-1,0,-1,1,0,-1,0,-1,1,2,1,1,-1,1,0,0,2,-1,0,0,1,0,0,2,-1,2,-1,-1,-2,0,1,0,1,1,0,0,2,1,0,1,0,2,1,0,1,-1,1,0,0,1,1,-1,1,0,-1,0,0,0,1,0,0,-1,-1,-1,-2,-2,2,2,0,0,-1,0,1,2,-1,0,1,1};
			57: counter1_out = '{-1,0,2,0,2,-2,-1,0,-1,0,0,-1,1,0,0,-1,0,1,0,1,-1,0,0,0,-1,-1,-2,0,0,0,-1,1,0,0,-2,-1,-2,-1,1,0,1,1,1,1,0,-1,-1,1,1,0,-1,-1,1,-1,0,1,2,2,2,0,2,1,0,0,1,0,-2,1,0,0,0,2,1,-1,0,0,0,2,-1,1,1,0,-1,1,-1,0,0,0,-1,-1,2,-1,0,-2,2,-1,-1,0,0,2};
			58: counter1_out = '{0,0,1,0,0,0,-1,1,0,0,2,3,-1,0,0,0,1,0,1,2,1,-1,0,-1,0,0,1,1,0,1,-1,0,0,-1,-1,-1,-1,0,0,0,1,-1,-1,0,0,-1,1,0,1,-1,-1,0,-2,1,0,2,-1,-3,2,2,0,-1,-1,2,-1,-1,-1,-1,1,1,-1,0,0,1,-1,2,0,0,-2,-1,0,1,0,-1,-1,-1,0,-1,2,0,0,2,-1,0,1,1,0,-1,-1,1};
			59: counter1_out = '{0,-1,1,2,-2,0,0,0,1,1,-1,0,-1,1,0,1,2,0,1,2,1,0,-1,2,-1,-1,0,-1,0,-1,2,0,0,0,-1,-1,-1,0,2,-1,-1,1,-1,-1,1,-1,-1,-2,2,-1,1,-1,0,-1,0,1,-1,0,0,1,2,0,0,-2,0,0,1,-1,-2,0,0,1,-2,1,1,-1,1,0,1,2,1,-1,0,0,0,0,-2,1,0,-1,1,0,1,1,-1,0,-1,1,2,1};
			60: counter1_out = '{1,0,0,0,0,1,-2,0,1,0,-1,-2,0,-1,-1,0,-1,0,1,2,1,0,2,-1,0,1,0,-1,-1,0,0,-1,0,0,0,0,0,-2,1,0,-1,0,2,1,-1,-2,-1,0,0,-1,-1,1,1,0,0,2,-1,0,1,0,3,2,1,0,-1,0,1,0,0,-2,-1,1,-1,0,-1,-1,0,0,0,0,1,1,0,1,-1,0,-1,2,-1,-2,1,0,-1,0,0,1,-1,0,0,0};
			61: counter1_out = '{0,1,0,-1,0,1,1,0,1,0,-1,0,-2,-1,0,-1,1,0,0,1,-1,0,0,3,1,-1,0,1,0,-1,0,0,-1,0,1,-1,0,0,0,-1,-1,-2,0,0,1,-2,1,-1,0,0,0,0,-1,1,2,0,1,0,-1,1,1,0,0,0,1,0,2,0,1,-1,0,2,0,0,1,1,1,-1,1,1,0,1,-2,-1,0,0,-2,0,0,-1,2,0,-1,2,0,1,-1,0,0,1};
			62: counter1_out = '{0,0,0,-1,-1,1,2,0,1,1,0,0,1,2,0,-1,1,0,-1,-1,-2,1,0,0,1,3,1,0,-1,0,1,0,1,-1,0,1,1,0,0,-1,1,1,-1,0,-2,1,0,0,0,2,0,0,0,0,0,0,-1,-1,-1,0,-1,-1,0,0,0,0,2,1,0,0,0,0,-2,1,1,-1,-1,1,1,-1,0,1,1,0,-1,0,0,-1,0,0,1,0,1,-1,0,1,0,3,0,1};
			63: counter1_out = '{1,1,-1,0,-2,-1,-1,0,0,1,1,0,0,0,0,-1,0,0,-2,0,0,-2,0,-2,0,1,-1,0,0,-2,0,1,1,0,0,-1,1,-2,1,0,0,1,0,-1,1,-1,-1,2,1,0,0,-1,0,0,0,-1,-1,0,-2,0,-1,-1,1,1,0,-1,1,-2,0,-1,0,-1,-1,1,1,-1,1,0,0,0,0,0,-1,1,-1,-1,-1,0,-1,1,1,2,-1,0,-1,-1,0,0,0,-1};
			64: counter1_out = '{0,-1,0,1,1,2,0,0,0,0,1,3,0,-1,0,-2,0,0,0,2,0,2,-1,1,1,0,2,0,0,0,-1,1,-1,1,-1,1,0,-1,-1,1,1,0,0,-1,1,-2,1,0,0,2,1,-1,0,1,-2,0,-2,1,-1,1,1,1,0,0,1,1,1,-1,-1,2,0,1,1,1,-1,0,-1,0,0,0,0,-1,1,2,-1,0,0,-1,1,0,1,1,2,0,0,0,-1,2,0,1};
			65: counter1_out = '{-1,0,0,0,0,-1,0,0,0,-2,2,-1,3,0,-1,1,-1,-2,-1,2,0,0,0,-2,-1,1,0,-1,1,0,2,0,1,0,1,0,2,0,1,0,2,-2,1,0,0,0,-1,1,-1,-1,0,1,1,0,0,-1,0,1,0,0,0,0,-1,2,1,0,0,0,1,-1,1,1,1,0,1,1,-1,-1,-1,2,2,1,2,0,0,0,1,0,-1,1,0,0,1,-1,-1,-1,-2,1,-1,0};
			66: counter1_out = '{0,-3,0,0,1,-1,0,-2,1,-1,-1,0,0,0,-1,0,0,0,0,-2,-1,1,-1,1,1,1,0,-2,1,1,2,-1,-1,0,3,0,0,-2,1,1,0,1,1,0,0,0,0,0,-2,-1,0,1,0,0,0,0,0,0,-1,0,1,-1,1,-1,0,0,0,0,0,0,1,-1,-1,-1,0,0,-1,0,0,-1,0,0,-2,0,0,1,-1,0,-2,-1,0,-1,0,1,-1,0,-1,-2,1,0};
			67: counter1_out = '{-1,-1,1,2,0,1,1,0,0,-2,0,-1,0,2,-1,-1,-1,-1,0,0,-2,0,1,-1,1,1,-1,0,-2,-1,0,1,0,0,1,-2,0,0,1,0,0,-1,0,0,-1,1,-2,-1,0,-1,0,0,2,1,0,0,-1,1,1,0,2,2,0,0,0,0,0,1,0,-2,-2,1,1,0,1,0,0,0,-1,0,3,-1,-1,0,2,-2,-2,0,0,-1,1,-1,1,1,0,1,-1,1,0,1};
			68: counter1_out = '{-1,0,1,3,0,-1,-1,0,-2,-1,1,0,-1,0,0,0,-2,0,0,-1,0,0,1,1,0,1,0,1,0,-2,1,-1,1,0,1,0,0,1,1,1,1,-2,0,2,0,1,0,-2,-1,-2,2,-2,-1,2,0,1,0,0,-2,0,-1,2,0,0,0,0,-1,0,0,0,1,0,-1,2,0,-1,-1,0,-1,0,1,0,-1,0,2,-1,0,-1,-1,0,1,0,2,0,1,-1,1,2,0,2};
			69: counter1_out = '{-1,0,2,1,1,2,-1,0,-2,1,-2,2,-1,1,-1,0,0,1,1,-1,-1,-1,-2,-1,0,-3,0,0,0,0,-1,-1,1,-2,-1,3,-1,0,0,-1,0,2,0,-2,-1,0,1,-1,1,0,1,2,0,1,2,0,0,0,1,-2,-1,-1,-3,1,2,0,0,1,1,1,-1,-2,-1,1,1,-3,-1,0,0,0,1,1,0,-1,0,0,-1,0,0,-1,0,0,-1,0,-1,1,0,0,0,1};
			70: counter1_out = '{0,-1,-1,1,1,2,2,-1,2,-1,-1,0,0,-2,-1,1,0,1,0,2,0,0,2,0,1,1,0,-1,-1,0,0,0,0,0,-1,0,1,0,0,-1,-1,0,0,0,0,2,0,1,-3,-1,0,0,-1,1,-1,-3,-1,-1,-2,0,-1,0,-1,1,-2,-1,0,0,1,0,0,3,-1,1,0,1,0,0,0,-1,1,1,0,1,2,-1,-2,1,1,1,-1,0,1,-1,0,2,-2,0,1,2};
			71: counter1_out = '{-2,1,-1,1,-1,1,0,1,-1,0,-2,-1,0,1,1,0,0,0,1,-2,1,0,0,0,0,-1,0,0,0,2,0,0,0,0,1,1,0,-2,0,-1,0,0,1,-1,1,-1,-1,1,-1,1,2,1,1,0,-2,-2,1,1,0,-1,0,0,0,0,0,-1,1,2,0,-1,0,2,-1,1,-1,0,0,-1,-2,0,0,1,-1,2,0,-1,-1,0,-1,0,-1,0,-2,-1,-1,0,2,-2,-1,-2};
			72: counter1_out = '{1,-1,1,-1,1,1,0,0,-2,-1,0,1,-1,-1,-2,-2,1,2,0,1,-2,1,-1,-1,0,-2,0,0,0,0,-1,1,0,2,1,1,0,0,0,1,0,0,1,0,-1,0,0,0,1,0,0,0,1,-2,0,-1,-1,0,-2,-1,2,-2,-1,1,-1,2,0,-1,1,1,0,1,0,1,-1,-2,-1,-1,0,0,-1,-2,-2,0,2,0,-1,1,3,1,0,-1,-2,0,1,1,-2,0,0,1};
			73: counter1_out = '{1,0,0,-1,1,1,-2,1,-1,0,2,1,0,1,0,-2,-1,0,1,1,1,-1,-1,-2,0,-1,1,0,-2,-1,-2,1,0,1,0,2,-1,2,2,1,-1,1,2,2,0,0,-1,0,1,0,-1,-1,-1,0,1,-1,2,1,-1,1,0,1,0,0,0,0,0,-1,0,-1,1,0,-2,-1,2,1,1,0,1,1,0,1,1,0,0,1,-1,1,0,0,0,-3,-1,-1,1,-1,-1,1,-1,2};
			74: counter1_out = '{0,0,0,1,0,-2,2,0,1,-1,2,-1,0,0,1,0,-1,0,0,0,0,0,0,-1,0,1,0,0,0,0,-1,0,-1,0,0,-1,1,0,1,2,-1,-1,0,1,2,-1,0,1,2,-1,-1,0,0,2,0,-1,0,1,-1,-1,0,1,0,2,0,-1,-1,-1,1,3,0,1,0,1,0,0,1,-1,1,-1,-1,1,-1,1,-1,1,-1,0,0,-2,0,1,-1,0,1,0,0,-1,-1,-1};
			75: counter1_out = '{1,0,1,-2,0,0,2,1,0,0,0,1,-2,0,-1,1,0,-1,-1,0,-2,0,-1,-1,1,-1,1,0,-1,0,-1,1,1,-1,-1,3,0,0,0,1,2,-1,0,0,2,0,1,-1,-1,-1,0,2,1,0,1,-1,-1,2,0,0,0,1,1,-2,0,0,2,-1,0,-2,0,1,0,1,0,0,0,-1,1,0,-2,-2,0,-1,-1,1,-1,2,0,0,1,1,0,0,-1,0,0,0,3,1};
			76: counter1_out = '{-1,1,0,1,-2,1,-1,0,1,0,1,1,-1,1,1,-2,-1,1,1,1,1,-1,-1,0,-1,-1,-2,-1,-1,-1,0,-1,2,1,-2,1,1,0,0,2,-2,-1,1,0,0,-1,-1,1,0,0,1,0,-2,0,1,0,0,-1,1,-1,1,0,-1,-1,1,0,1,-1,1,0,1,1,-1,0,-1,0,1,0,0,0,-1,2,1,2,-1,1,2,0,-1,-1,0,0,0,0,-1,0,-2,-1,0,0};
			77: counter1_out = '{-1,0,0,1,-1,1,1,1,0,0,1,0,-1,1,0,0,-1,1,-1,0,-1,-1,-1,-1,-2,1,-1,2,-1,-1,-2,1,0,-2,0,1,-2,-1,0,2,0,0,-2,0,0,0,-1,1,0,-1,-1,-1,2,0,0,2,-1,2,-2,0,0,0,0,1,-1,1,0,0,0,-1,-1,0,1,-1,1,0,0,1,-1,1,-1,1,-1,0,0,2,2,-1,0,2,-1,0,0,0,-1,2,-1,1,1,0};
			78: counter1_out = '{0,-1,0,0,0,0,-1,1,0,-1,0,0,-1,0,-1,0,-2,0,1,2,1,1,0,-2,0,0,1,-1,0,-1,1,-2,0,0,1,1,1,-1,2,0,1,-1,0,-1,0,1,2,-1,-1,-2,1,-1,1,-1,0,1,1,-1,0,0,2,1,0,2,0,-1,1,0,2,-2,-1,0,-1,0,0,-1,0,-1,-1,-1,-3,0,-1,-1,-3,0,0,1,0,2,0,1,0,0,1,1,1,0,-1,-1};
			79: counter1_out = '{0,1,1,-1,1,-1,0,-1,3,1,1,0,2,0,1,0,0,0,0,0,0,2,-2,2,1,0,-1,-1,-1,-1,-1,2,1,1,0,1,0,2,-1,0,-1,0,2,2,1,-2,1,0,-2,-1,0,0,-1,0,0,0,0,-1,-3,1,0,-1,2,1,-1,-1,0,-1,1,0,1,1,0,0,-1,1,-1,-2,1,0,-1,0,-1,1,0,-1,1,0,2,1,0,-1,0,1,-2,1,1,-1,0,2};
			80: counter1_out = '{1,-2,-1,0,-1,-2,0,-2,0,0,-1,0,-1,-2,0,-1,0,1,1,0,-1,1,2,1,1,-1,0,1,0,1,0,-1,0,-1,0,1,-1,0,1,2,-2,1,0,1,1,0,0,1,-1,0,0,0,1,-1,-1,-1,1,-1,1,-1,-1,1,0,0,-1,1,-1,0,0,1,0,-1,0,0,1,1,0,3,1,0,0,1,0,1,0,0,1,0,-1,-1,1,0,0,-1,-2,-1,-1,0,1,0};
			81: counter1_out = '{1,-1,2,0,-2,0,1,-2,-1,0,-2,2,1,1,-1,0,0,0,0,-1,-1,-1,-1,0,2,-1,-2,1,-2,-1,-1,0,1,1,0,0,1,0,0,0,0,1,0,1,0,0,0,1,1,0,2,0,-1,2,-1,2,1,0,-1,-1,-1,0,-1,0,0,1,-1,-1,0,-1,1,1,-2,-1,0,-1,0,0,0,0,1,-1,0,0,2,-1,-1,-1,1,0,0,0,1,0,-2,0,-2,1,0,1};
			82: counter1_out = '{0,-1,1,-1,-1,0,-1,2,2,0,0,0,1,1,0,-1,1,-1,1,1,1,0,1,0,-1,1,0,0,0,-1,-1,1,0,1,-1,-1,0,1,0,1,0,0,0,1,0,1,2,2,0,0,0,1,1,-2,1,0,0,1,0,0,2,0,2,2,0,0,1,0,-2,1,-1,0,1,-1,-1,2,-1,2,2,-1,-1,-1,-1,-1,-1,0,0,-2,-1,1,-1,-1,1,0,1,0,1,1,1,0};
			83: counter1_out = '{-1,0,-1,2,-1,0,0,1,0,0,-1,3,-1,0,0,2,0,0,-1,0,-1,1,0,1,1,0,0,-1,1,0,-1,0,0,0,0,1,-1,2,-2,-2,-1,-1,-2,1,1,0,2,0,-2,0,-1,1,0,0,-1,-2,-1,1,1,0,1,-1,-1,-1,0,1,-2,1,-1,2,-1,-1,-1,0,0,0,1,1,1,2,1,1,0,0,0,0,-1,1,1,1,-1,0,-1,2,-1,-1,1,1,0,-2};
			84: counter1_out = '{-1,-1,-2,1,-1,0,0,0,1,2,-1,1,0,-1,0,0,0,-1,-1,-1,-1,-1,0,-1,1,-1,0,2,1,0,-1,-1,0,-1,1,0,2,1,0,1,-2,-1,-2,0,-1,1,0,1,-1,1,2,-1,0,2,0,-1,1,1,-1,1,0,-1,-1,-1,-2,0,-2,1,1,0,0,-1,2,0,1,1,0,0,1,-1,0,0,-1,0,-1,-1,1,0,1,0,1,1,1,-1,0,-1,0,-1,-1,1};
			85: counter1_out = '{0,-1,1,1,-1,0,-1,-1,0,0,0,1,0,1,-1,-1,1,-1,1,-1,0,-2,-1,0,0,0,0,-1,-2,-1,1,0,-1,0,0,-2,1,-1,0,0,0,1,0,-1,-1,0,-1,0,1,-1,0,-2,-1,0,-2,0,0,2,0,0,0,0,0,1,-1,0,-2,1,0,0,0,0,1,0,-1,1,1,0,0,-2,-1,0,1,-1,-1,0,-1,0,-1,-1,0,1,-1,0,0,1,2,1,1,0};
			86: counter1_out = '{-2,0,1,1,0,1,-1,1,1,0,-1,-2,-1,0,1,2,-1,-1,1,-1,1,0,1,-1,0,-1,-1,0,1,-1,-1,0,0,0,-2,1,2,0,1,-2,-1,2,0,-1,0,0,-1,0,0,2,1,0,1,0,0,0,1,-1,1,1,-1,0,0,-2,1,1,-2,0,0,-2,-1,0,2,0,0,1,0,-1,2,-1,-1,0,-1,0,-2,1,0,0,-1,-1,1,0,-2,-1,2,-1,-1,2,1,1};
			87: counter1_out = '{0,1,1,0,0,-1,0,0,-1,-1,0,1,1,-1,-1,-1,-1,0,-1,1,2,0,1,-1,0,0,-1,1,0,1,0,2,0,0,0,2,0,0,0,1,2,1,1,1,2,1,-1,0,1,-2,0,-1,-1,-1,1,0,-1,1,-1,1,0,1,1,1,-1,0,-1,-1,2,-1,1,0,0,0,-1,-1,1,1,-1,1,2,2,-1,-1,0,-1,0,-1,-1,-1,1,0,-2,0,1,0,0,0,0,0};
			88: counter1_out = '{0,0,0,1,1,0,0,0,1,-1,0,0,0,2,-2,1,1,2,0,0,1,-1,0,-1,-1,-2,0,0,0,-1,0,-3,0,1,0,0,0,2,-1,0,0,0,0,0,-1,0,1,1,-1,3,1,0,-1,-1,-1,0,1,1,1,1,0,1,-3,-1,-1,1,0,2,0,0,-1,-1,0,2,0,2,0,0,1,1,-1,1,0,0,-2,0,0,0,0,1,-1,0,-1,-1,1,1,0,-3,0,-1};
			89: counter1_out = '{0,2,1,2,1,0,1,0,1,-1,-1,-1,1,-2,1,1,1,2,1,1,1,2,0,-1,-2,-1,-2,-1,0,0,-1,-1,-1,-1,-1,0,1,-2,1,-2,-1,0,0,-1,-1,2,0,-1,0,0,0,1,-2,-1,-1,1,0,0,0,2,0,0,0,0,1,-1,0,-1,0,0,0,1,1,1,0,-1,1,0,1,-2,1,1,-1,1,2,-1,2,0,0,-1,1,0,-1,-1,1,1,1,-1,-3,0};
			90: counter1_out = '{-1,-1,1,1,-1,0,1,-2,-2,-1,1,-1,-1,1,1,0,1,0,0,-1,-1,0,1,-1,-1,0,0,1,1,2,0,0,1,1,1,0,0,0,1,1,-1,1,-1,-2,2,0,-1,-1,0,1,0,-1,1,2,0,-1,1,0,0,1,0,-1,0,-1,-1,0,-1,-1,0,0,-1,-3,0,1,-1,1,1,-1,-2,1,0,0,0,1,0,0,-1,-2,0,1,1,1,0,0,-1,-1,-2,-1,0,0};
			91: counter1_out = '{1,-2,0,1,1,2,0,-1,0,0,0,1,-1,2,-1,1,2,0,0,0,-1,1,0,0,0,1,1,-1,1,1,-2,0,1,-1,-1,2,0,-1,0,-1,1,-1,-1,1,-1,1,-1,-2,0,0,-2,0,0,0,0,-1,0,1,-2,0,-2,0,3,0,0,-2,0,1,0,1,1,0,-1,0,-1,-1,0,1,0,-1,-2,0,0,-1,1,-1,0,3,1,1,1,1,-3,3,0,-1,0,0,2,-1};
			92: counter1_out = '{1,0,1,1,0,-2,1,-1,0,0,-1,0,0,0,1,0,-1,-1,1,0,0,1,-2,-2,1,0,1,-1,0,0,-1,0,0,-1,0,-1,2,0,0,-1,0,-1,0,0,-1,0,-1,1,0,0,1,1,0,0,1,0,0,-1,-1,0,1,-1,1,0,1,0,-1,0,0,2,-2,0,1,0,0,-1,0,-1,0,0,0,0,2,-1,0,0,-2,-2,2,-1,-1,0,-2,1,0,0,-1,0,0,0};
			93: counter1_out = '{-2,0,1,2,1,0,-1,-1,-1,1,1,0,1,0,0,1,0,0,0,-1,-2,0,0,0,0,-2,1,-1,0,-1,-1,-1,2,0,0,0,-1,2,0,-1,1,0,1,1,-1,1,-1,0,1,2,0,-1,1,0,-2,1,-1,1,-2,0,1,1,-1,-1,0,0,-1,0,-1,0,0,0,0,0,0,-1,1,0,-1,0,-2,0,-1,-2,-1,1,-1,-2,-1,0,0,-2,0,0,1,0,1,-2,-1,0};
			94: counter1_out = '{0,1,0,0,1,0,1,1,-2,2,-1,1,0,1,1,0,1,0,-2,2,0,-1,-1,0,1,2,0,1,-1,1,0,2,0,-2,0,1,1,-1,0,0,-1,0,0,0,0,0,-2,1,0,1,0,0,-1,1,1,1,1,0,-1,-1,1,0,-1,1,0,1,-2,2,1,-2,0,-1,1,-1,2,-1,-3,0,0,0,0,0,3,1,1,-1,0,1,1,-1,1,-1,1,0,1,0,1,0,0,-1};
			95: counter1_out = '{1,1,2,0,0,0,4,-1,2,0,0,2,-1,0,-1,-1,0,0,-1,-2,1,0,0,-1,1,1,0,1,-1,-1,0,2,0,2,0,0,-1,-2,0,1,-1,2,1,0,1,-1,0,0,-2,1,0,2,-1,-1,-1,-1,-1,-2,0,-2,0,-1,-1,0,1,0,1,0,-1,-1,-1,2,-1,-1,0,0,-2,0,-1,-1,0,0,-1,0,0,1,-1,-1,-1,0,1,0,0,-2,0,1,1,0,1,1};
			96: counter1_out = '{-2,1,-1,1,0,1,-1,-2,-1,-1,1,0,0,1,-1,-1,1,1,0,0,-2,-1,1,1,2,-1,2,-1,-1,0,0,-1,0,1,-1,1,0,0,1,-1,1,0,0,-1,-1,-1,-1,0,0,2,0,0,0,2,0,0,-1,-1,-1,0,4,0,0,0,0,-1,-2,1,0,-1,1,0,1,0,0,-2,1,-2,0,-2,1,1,0,-1,0,0,-1,-2,0,0,-2,-2,2,1,0,-1,-1,0,0,0};
			97: counter1_out = '{0,1,0,-1,1,-2,3,-1,-1,0,-1,0,1,0,0,0,1,2,1,1,0,0,1,0,1,-1,0,0,-2,-1,1,-3,0,0,1,0,0,0,0,-2,1,0,1,0,1,0,1,0,0,0,1,0,-1,0,-1,-1,0,-1,-1,0,-1,-1,-2,0,0,1,0,1,1,-1,1,1,-2,2,2,1,2,1,0,-1,0,1,0,0,1,-2,0,-3,1,0,-2,0,1,1,-1,-1,2,-1,-1,1};
			98: counter1_out = '{-1,0,0,0,1,1,-1,1,0,-1,0,0,2,1,-1,-1,0,-1,1,1,-2,-2,0,0,-1,0,0,0,0,2,1,1,0,0,-1,1,2,2,2,-1,0,-2,0,0,-1,0,-1,1,1,1,1,0,0,0,1,0,0,0,-2,0,2,2,0,0,-1,1,1,1,1,-1,1,-1,1,0,1,1,-2,-1,1,-1,0,-1,-1,-2,1,-2,0,-1,0,0,1,-1,-2,-1,1,1,1,-1,-1,0};
			99: counter1_out = '{0,-2,1,0,0,-1,-2,0,0,-1,1,0,0,-1,1,0,-2,0,-2,0,0,-1,0,-2,1,-1,1,-1,-2,-1,2,1,-1,1,1,-1,2,0,-1,0,2,0,1,1,1,0,0,0,-1,2,0,2,0,2,-1,1,-2,2,-1,0,0,1,-3,2,1,-1,-1,1,0,1,0,-3,-1,0,0,-2,0,-1,1,0,1,0,0,0,0,0,0,-1,2,0,0,1,0,1,2,0,0,0,2,-1};
			100: counter1_out = '{0,0,0,-2,-1,1,-1,0,0,-2,0,3,0,0,0,2,0,-1,-1,0,-1,-1,1,0,0,2,1,1,-1,1,0,0,-1,-1,1,-1,0,0,1,-2,0,-3,0,0,0,0,0,0,-2,0,-1,1,2,1,-1,0,1,2,-3,0,0,0,1,0,0,1,-1,-1,-1,2,0,0,0,-1,0,1,-2,0,1,0,-2,0,1,0,0,1,0,0,0,0,0,-2,-1,1,-2,0,2,1,0,-1};
			101: counter1_out = '{-1,0,2,-1,0,1,0,1,2,-2,-1,-1,-1,0,0,-1,-1,0,0,0,1,0,0,-1,0,0,1,0,0,0,0,-1,-2,-1,0,0,0,0,0,-1,0,0,1,0,-1,1,-1,-2,-1,0,0,-1,0,-2,-1,1,0,-1,-2,-1,2,1,-1,0,1,-3,2,1,-1,3,0,0,-1,0,0,4,0,0,1,1,1,-1,1,0,2,0,0,1,-1,0,-3,0,0,0,0,0,2,1,0,0};
			102: counter1_out = '{0,0,3,0,-2,-1,0,0,-1,-1,-1,1,0,0,0,-1,1,1,-2,0,0,-2,0,0,-1,1,0,0,0,0,1,1,-1,0,2,1,-2,-1,1,-1,1,-1,1,-1,1,2,0,0,-1,-1,0,0,1,-2,-1,-2,-1,1,-1,0,0,2,0,0,-1,1,0,1,2,-1,1,1,0,-1,1,1,1,-1,1,-1,0,0,0,0,0,0,-1,0,0,0,1,-1,1,1,-1,1,0,0,-1,-1};
			103: counter1_out = '{1,-1,0,-1,0,1,-2,-2,1,1,-2,1,-1,-2,-1,-2,0,0,0,1,0,0,0,1,-2,1,1,0,-1,0,1,1,0,0,0,1,0,0,0,-1,0,1,0,-1,-1,-1,1,1,-1,-1,-1,0,0,1,0,0,1,1,-1,1,1,-1,-1,0,-1,1,-2,1,0,1,0,0,-1,-1,-1,1,0,0,2,0,-1,-1,-2,0,1,1,0,0,0,2,1,-1,0,-1,0,1,0,0,1,0};
			104: counter1_out = '{1,1,2,-1,1,1,1,3,1,1,-1,0,0,1,0,1,-2,0,0,0,0,-2,0,-1,0,0,-1,-1,2,-2,-1,-2,0,0,0,0,-1,1,1,0,0,-1,1,0,0,1,-1,2,-1,0,1,-2,1,1,0,-1,1,2,1,-2,0,-1,0,-2,2,-2,0,0,2,-1,1,1,-1,0,2,-1,0,1,0,0,0,-1,-2,1,1,1,1,1,1,-1,-1,1,-1,0,-1,1,0,2,1,1};
			105: counter1_out = '{0,1,1,1,0,0,-1,-1,1,0,0,-2,1,1,-1,1,1,1,-1,0,-1,-1,0,0,1,1,-2,0,-3,1,1,0,-1,0,2,1,-1,1,0,0,1,-2,0,2,1,-1,0,-1,0,-1,-1,0,1,1,-1,-1,0,1,-3,2,0,0,0,1,0,1,-3,-2,-1,1,-1,-2,1,-2,-1,1,0,1,-1,0,0,-1,-1,0,-2,0,-1,1,1,1,-1,0,0,-1,1,0,-1,1,0,-1};
			106: counter1_out = '{2,-2,0,-1,-1,0,0,-1,0,0,0,0,1,-1,-1,2,-1,0,0,0,1,0,-1,2,-1,0,1,1,0,0,0,1,-1,1,-1,-2,2,0,0,0,-1,-1,-1,1,0,0,1,0,1,-2,-1,1,1,-1,0,-1,-1,2,0,1,0,0,-1,-2,-1,1,1,0,0,0,-1,-1,0,1,-2,0,-1,2,0,0,0,-1,1,-1,0,-3,1,2,-1,2,1,-1,-1,1,1,0,1,-2,0,0};
			107: counter1_out = '{0,-1,0,-1,0,0,1,0,1,1,0,-2,0,3,0,0,0,0,1,0,0,1,0,-1,0,-2,1,0,-1,-1,-1,-1,-1,-1,0,-2,0,-2,1,1,0,0,2,2,-1,1,0,0,-1,-1,0,-1,0,0,1,-2,-1,-1,0,1,-1,0,1,1,1,2,1,0,2,-1,-2,0,1,1,0,-2,1,-2,1,0,-2,0,-1,-2,2,2,1,0,1,1,1,0,2,1,1,1,0,1,1,0};
			108: counter1_out = '{0,-1,0,-2,1,0,-1,-1,2,0,0,0,0,-1,-1,-1,1,-1,1,-1,0,0,1,1,0,-3,1,-1,1,1,-1,-1,0,0,0,-2,-1,-2,-1,1,1,-1,0,1,0,1,-2,-1,0,1,0,1,1,0,1,1,-1,0,-1,0,0,2,2,-3,-1,0,0,-2,-1,-1,1,0,0,0,0,0,-1,0,0,1,2,1,1,0,1,-1,1,0,1,1,-1,1,0,0,0,0,1,1,1,0};
			109: counter1_out = '{0,0,0,-2,0,0,0,1,0,1,1,0,0,1,-1,-1,0,-1,0,1,0,0,0,2,2,0,0,1,0,1,-1,0,0,2,-1,0,-1,-2,1,-1,0,1,0,-1,1,0,1,-1,-1,0,1,1,1,1,-1,0,0,0,-1,1,1,1,-1,1,-1,0,0,0,-2,0,2,-1,-2,0,0,0,1,0,0,1,0,0,-2,0,-1,1,0,0,0,0,0,2,-3,-1,1,0,0,1,1,0};
			110: counter1_out = '{0,-1,-1,1,-1,0,1,0,-1,-2,-1,1,-1,0,0,0,0,-1,0,-1,1,1,1,0,1,0,2,0,0,-1,-1,-1,1,-2,1,1,-1,-3,1,-1,-1,-3,-1,1,1,-2,1,-2,1,1,-1,1,0,-1,1,2,-1,-1,0,0,-1,0,-1,0,0,0,1,0,-1,0,1,0,0,0,-1,0,-1,1,-1,2,0,-2,1,0,1,-1,1,-1,-1,2,0,0,0,2,0,-1,0,2,2,1};
			111: counter1_out = '{1,0,2,0,-1,-1,0,0,1,-1,1,1,1,-1,0,-1,0,1,0,-2,-1,0,-1,-1,0,0,0,-1,2,-1,2,0,-1,0,-1,-1,-2,-1,-1,2,-1,-1,1,1,1,0,0,-1,1,1,0,1,0,0,1,1,0,-1,0,0,-1,0,1,0,0,0,1,0,-1,-1,2,0,1,0,1,-3,-1,-1,2,0,1,0,-2,1,0,0,-1,-1,-1,-2,0,1,2,-1,1,1,2,0,-1,-1};
			112: counter1_out = '{1,0,-1,1,0,0,0,0,2,0,0,2,0,0,0,0,-1,-2,1,2,-1,-1,1,0,0,-1,1,0,0,-1,1,-2,0,-1,0,2,1,0,-2,0,1,-1,1,-1,0,0,1,1,1,0,0,-2,0,1,0,0,-1,-1,0,1,0,0,0,0,0,1,0,2,-1,0,2,-1,0,0,1,1,1,0,0,0,0,0,-1,-1,0,-1,-1,0,1,0,0,0,0,1,0,-1,-2,1,0,-3};
			113: counter1_out = '{-1,0,1,0,1,-2,-1,-1,-1,1,-1,2,0,1,-1,1,0,1,0,0,0,1,1,-1,-1,-1,1,0,1,-1,1,-1,2,0,0,1,0,1,2,0,0,1,-2,-2,0,-1,-1,-1,1,-1,-2,0,-1,0,1,2,-2,-2,1,2,1,0,-3,-1,0,0,-1,0,1,1,-1,2,1,0,1,1,2,-1,-1,1,-1,0,-1,0,1,2,1,0,-1,-1,0,-1,-1,1,0,0,0,-2,1,0};
			114: counter1_out = '{0,2,-1,0,0,1,-3,0,0,0,0,1,0,-1,0,-1,0,0,0,0,1,0,3,1,1,-1,1,1,0,0,2,0,0,0,0,1,0,-2,0,0,1,-2,0,1,-1,1,-1,0,0,-1,0,1,1,-1,-2,0,0,1,-1,-1,-1,1,-1,-1,-3,2,0,1,-2,-1,0,-1,2,1,0,1,1,-1,-1,1,0,0,0,2,0,0,2,0,0,1,0,-1,-1,-1,-1,-1,1,0,0,0};
			115: counter1_out = '{-2,2,0,0,0,-2,0,1,-2,1,0,0,2,0,0,-1,-2,-1,0,0,-2,-1,0,0,0,2,0,-1,0,-1,0,0,-1,1,1,2,1,1,0,1,1,0,-1,0,1,-1,2,1,2,0,0,1,-1,1,-2,0,1,-1,-1,1,1,1,-2,-2,-1,1,-1,-1,0,1,-3,-1,1,-1,0,1,0,0,0,0,0,-1,1,1,-1,-2,-1,0,-1,0,1,-1,0,1,-1,1,-3,2,2,-1};
			116: counter1_out = '{-1,0,-1,-1,1,2,-1,0,-1,1,1,-2,1,-1,0,-1,-1,-1,-1,1,-1,-1,-2,-2,-1,0,1,-2,0,0,-1,1,-1,0,-1,2,2,1,0,-1,1,0,-2,-1,-1,0,1,0,-1,-1,0,1,1,1,0,1,0,-2,0,0,-1,0,-1,-2,1,-2,-1,-2,0,-2,-1,1,0,1,1,0,1,-1,0,0,-1,0,-1,0,1,1,1,-2,0,1,-3,0,1,0,0,-1,-2,1,2,0};
			117: counter1_out = '{1,0,0,2,0,0,1,-2,0,1,0,-1,0,2,1,-1,0,0,0,-1,-1,0,0,0,1,0,1,1,0,0,0,1,0,1,1,0,0,0,-3,-2,1,0,-1,0,0,0,0,2,-1,0,1,-1,1,-1,0,0,-2,0,0,-2,1,-1,0,0,1,1,-1,-1,0,0,-1,-2,0,-1,0,1,-1,1,0,2,0,1,0,1,0,0,-2,-1,-2,-1,0,0,0,0,-1,-1,-1,0,-1,0};
			118: counter1_out = '{-1,0,2,1,0,2,0,2,-1,0,0,-3,1,1,-1,0,-2,1,0,0,0,0,-1,0,1,1,1,0,-1,0,0,0,1,0,-1,2,0,1,0,-1,0,2,1,-1,1,-1,0,1,2,1,-1,0,1,1,2,-1,-1,-1,0,0,1,1,-1,0,0,0,-1,0,0,1,1,-1,-1,0,0,0,2,1,-1,0,1,0,1,-1,-1,0,0,-1,1,-1,-1,2,1,-1,0,-1,1,1,1,-2};
			119: counter1_out = '{1,0,0,1,1,-2,-1,-1,0,0,-1,1,-2,-1,1,1,1,1,1,1,1,1,0,-1,0,-2,0,0,1,1,0,0,0,0,0,0,-1,-1,0,0,0,0,0,1,0,-1,0,0,1,-1,0,-1,1,1,2,0,2,-1,0,1,1,2,3,1,1,1,-1,-1,-1,-2,0,-1,0,0,1,1,1,1,1,0,0,-1,0,1,2,1,-1,1,0,-1,0,1,0,-1,1,-1,0,0,-1,0};
			120: counter1_out = '{0,2,1,-2,-1,-1,-1,0,-1,0,0,-3,1,0,0,-1,1,-1,-2,-1,1,0,0,1,1,-1,0,-1,0,0,0,0,-1,1,1,-1,0,-1,0,2,0,0,-1,0,0,1,1,0,0,1,0,-1,-2,-1,1,-2,0,0,0,-1,1,-1,-1,0,-2,-1,0,1,0,1,1,1,0,0,0,-1,0,-1,0,-1,0,0,0,0,0,-1,0,-1,0,-1,1,1,0,1,-1,-1,2,0,0,-1};
			121: counter1_out = '{1,1,0,-1,-1,0,-1,1,1,0,0,0,0,-2,0,0,-1,-1,0,2,-1,-1,2,1,1,0,0,0,-1,1,1,0,2,-1,0,2,-2,1,1,0,0,0,-1,0,1,-2,2,0,-1,-1,1,-1,1,1,0,0,1,1,-1,-1,2,1,0,-1,1,1,0,0,0,0,-1,0,-2,1,2,-1,0,1,-1,1,-1,2,1,0,1,2,0,0,0,0,-1,0,-1,1,1,1,0,0,0,2};
			122: counter1_out = '{0,0,-1,0,1,0,-1,0,0,-1,0,0,-3,1,-1,-2,0,0,2,0,1,2,-1,0,-2,-1,1,0,0,-2,1,-1,0,1,0,0,0,0,1,0,-1,-2,2,-2,0,-2,-1,1,2,2,-1,-1,-1,0,-1,-1,-1,-1,-3,0,1,1,-2,0,0,1,0,-1,2,0,0,0,0,-2,0,0,1,1,2,0,-2,-2,0,1,1,-2,0,0,-1,0,0,0,1,1,0,-1,0,-1,-1,0};
			123: counter1_out = '{1,0,1,-2,0,-1,-1,0,1,1,0,-1,2,0,1,0,0,0,1,-1,0,1,1,-2,0,-1,-2,0,0,1,1,0,1,0,-1,1,1,-1,1,1,-1,1,1,-1,0,-1,0,0,1,0,1,-2,0,-1,0,-1,1,-1,-1,2,3,1,0,0,0,1,-2,0,3,0,-2,2,1,1,1,1,-1,0,-2,2,1,0,2,-2,-1,2,-1,-1,0,0,1,1,0,0,1,1,1,-1,0,0};
			124: counter1_out = '{1,-2,0,1,1,0,2,-2,2,1,0,0,1,0,0,0,1,0,-2,2,-2,0,0,0,0,0,0,-1,-1,0,0,0,-1,-1,1,-1,-1,-2,2,0,0,-1,2,0,-1,0,1,0,-1,2,0,0,0,0,1,0,0,1,-1,-1,0,1,0,-1,2,0,0,1,-1,-1,0,1,-1,1,1,-1,1,0,1,-3,0,1,0,0,0,-1,-2,1,0,0,-1,-1,0,0,-2,-1,2,1,0,-1};
			125: counter1_out = '{2,0,1,0,0,-1,1,1,1,-1,-1,2,-2,0,0,-1,1,0,0,-2,-1,1,0,0,-1,-2,2,0,-2,0,0,-1,-2,-1,2,0,1,-1,-1,3,1,-2,3,-2,-1,1,-1,-1,2,-1,1,0,0,-1,1,0,-2,-1,-2,0,1,0,-1,-1,0,1,-1,1,1,0,0,0,1,1,0,0,0,0,-1,2,0,0,0,0,0,-1,0,0,0,-1,0,-1,0,0,1,1,0,0,-1,2};
			126: counter1_out = '{-1,-1,-1,-1,2,-1,1,1,0,0,1,-1,0,1,-1,1,1,-2,-1,1,-2,0,1,-1,-1,0,1,0,0,0,1,-1,0,-2,1,-2,-1,-1,-2,0,0,1,2,1,0,-1,0,0,1,-1,0,0,0,0,0,0,1,0,-3,0,0,0,-2,-1,2,3,1,1,2,0,-2,-1,1,1,0,0,-1,1,0,2,2,0,0,2,0,-1,1,-1,1,-1,-1,-1,0,-1,0,2,0,0,2,0};
			127: counter1_out = '{1,0,-1,1,-1,0,2,2,0,0,-1,2,-1,-1,1,1,1,-1,-1,1,-1,0,1,-2,1,-1,1,0,0,0,-1,-1,1,-1,1,1,1,-2,0,1,1,-1,4,2,-1,0,-1,0,-1,0,2,0,0,-1,0,2,0,1,-1,1,-1,1,-1,0,0,0,2,-1,0,1,-2,-4,-2,-1,-2,0,1,0,1,1,1,0,0,1,0,-1,-1,-1,-1,1,2,0,-1,-1,1,1,3,1,0,-1};
			128: counter1_out = '{0,0,-2,0,0,0,0,-1,1,0,0,0,0,-1,-2,1,2,1,0,0,0,-1,0,2,0,0,1,1,-1,1,-1,0,1,1,3,1,2,0,1,1,1,0,0,0,0,-1,1,0,-1,1,0,-1,1,-1,-2,0,1,1,0,-1,-1,1,-2,-1,1,1,1,0,1,1,0,0,1,-1,1,-1,1,0,0,-1,0,0,1,1,-2,-1,-1,0,1,-2,-1,2,0,0,-2,0,1,-1,0,2};
			129: counter1_out = '{-1,1,-1,-1,0,-1,0,0,1,0,-1,1,0,-1,0,0,2,1,0,1,-1,0,1,0,0,0,1,1,-1,2,-1,0,1,1,0,0,1,0,1,0,0,-2,0,-1,1,1,-1,0,1,-1,-1,-1,0,0,1,0,0,0,2,2,-2,1,1,-1,1,0,2,0,0,-1,1,1,-2,3,1,-2,0,0,-1,0,3,0,-3,-1,-2,1,0,0,1,-1,-1,-1,0,0,0,0,0,1,0,2};
			130: counter1_out = '{-2,-1,1,0,-1,0,-1,1,0,2,-1,2,1,1,0,1,2,-2,1,1,0,-1,1,0,-2,1,0,0,0,1,-1,0,0,-1,0,0,1,1,1,0,1,0,-2,1,0,0,0,-1,0,2,1,-1,1,0,-1,-2,0,1,1,0,1,-1,-1,1,1,0,1,-1,2,-1,0,2,-3,0,-1,0,2,-1,2,2,1,-1,0,-1,0,-3,1,1,0,-2,0,0,-2,0,0,1,1,-1,-1,0};
			131: counter1_out = '{0,-2,-1,0,1,1,0,0,-1,0,0,-1,-1,0,1,2,0,0,0,-1,1,-1,-1,0,0,0,2,-1,-1,0,1,0,1,1,1,1,0,-2,1,0,0,0,1,1,1,1,0,-2,0,1,0,0,0,1,0,0,-1,0,-3,0,0,-1,-2,1,2,0,0,0,0,-1,1,0,0,0,1,0,2,-1,-1,0,-2,-2,0,0,0,0,-1,2,1,-1,-1,-1,0,0,-1,-1,1,0,-1,2};
			132: counter1_out = '{0,1,0,-1,-1,0,-1,-2,-2,0,1,1,0,0,1,-1,0,-1,-1,0,2,0,0,1,0,-1,-1,0,0,-2,0,0,1,0,1,-2,1,-1,0,0,2,1,1,1,-1,1,-1,-1,-3,-1,0,0,0,-1,-1,-1,-2,1,0,0,0,-1,0,0,-1,-1,1,-2,1,1,-1,1,0,-1,0,2,-1,1,0,1,-1,-3,-1,0,0,0,-2,2,-1,1,0,-1,0,1,1,2,0,0,-1,2};
			133: counter1_out = '{1,2,0,1,0,-1,2,0,-2,2,-2,-1,0,-1,-1,0,0,-1,1,-1,0,-1,0,0,-1,1,-1,0,2,-1,-1,0,0,2,-1,-1,-1,0,1,2,0,0,-1,2,1,-2,0,-1,1,0,0,-1,-1,0,0,1,0,0,0,1,1,0,-1,-1,0,0,0,1,0,1,0,-1,1,0,-2,-1,3,1,-2,-1,-1,0,-2,0,0,-1,1,0,0,-1,1,2,-3,0,1,1,-2,0,0,1};
			134: counter1_out = '{1,0,0,-1,0,-2,0,0,0,-1,-1,1,-1,-1,1,1,-2,1,0,0,1,-1,-1,-1,0,0,0,-1,0,0,0,-1,1,0,0,0,-1,-1,-1,0,0,-2,-1,1,1,1,-2,0,1,0,-1,0,0,0,1,-1,-1,-1,0,2,-1,0,-2,-1,1,0,-1,2,-1,-1,-1,-1,-1,-1,0,1,1,0,1,0,-1,0,-2,-3,-2,-2,-1,1,0,1,0,2,0,2,0,2,0,-1,1,-1};
			135: counter1_out = '{0,-1,-1,0,0,0,1,-1,2,1,-1,1,0,2,0,2,-1,1,0,0,2,0,0,1,0,2,-1,-1,0,-1,0,2,1,0,0,-2,1,1,-1,1,1,0,0,0,0,1,-1,0,-1,1,-1,0,0,-2,0,-1,2,1,0,0,0,0,1,-1,0,1,2,1,1,-1,0,1,1,2,-2,-2,0,0,1,0,0,-2,0,1,1,0,-1,1,0,0,-1,0,-1,1,-1,-2,-1,1,1,-2};
			136: counter1_out = '{0,0,0,-1,0,-2,0,-2,1,1,0,1,2,0,0,-1,0,-1,-2,0,1,0,0,0,1,0,0,-1,1,-1,-1,1,0,1,0,0,-1,-2,4,0,-1,1,0,1,-2,0,2,-2,0,-1,0,-2,0,1,-1,0,1,-1,1,-1,0,1,0,-1,0,1,1,0,1,1,-1,-1,1,1,-2,0,1,0,0,1,1,0,1,0,-1,0,0,1,1,-1,0,1,-1,0,0,-1,0,1,1,1};
			137: counter1_out = '{1,2,2,2,0,-1,-1,1,0,0,0,1,-1,0,-2,0,-2,0,-1,0,-2,1,-2,0,-1,-1,-1,0,0,-2,0,1,-1,-1,0,1,0,-1,1,-1,-1,-1,0,0,1,1,1,1,0,1,0,0,-1,1,-1,-1,-2,-2,0,0,-2,1,1,1,1,-1,0,0,0,0,1,1,1,1,1,0,-2,0,0,-1,-1,2,2,1,0,0,1,-1,0,1,0,-1,0,1,0,2,-1,0,2,0};
			138: counter1_out = '{-1,0,1,2,0,-1,0,0,-2,1,-2,-1,1,-1,1,0,1,-1,2,-1,0,-1,-1,0,-2,0,1,1,0,-1,1,0,2,2,-3,0,0,0,0,-1,-1,-1,0,-1,0,0,-1,0,-2,1,1,1,0,-1,-1,-1,-2,0,0,0,-1,0,1,1,0,0,0,0,-2,1,-2,1,0,0,1,-1,-2,0,1,0,0,1,0,-1,0,0,0,0,-1,-1,0,-1,1,-1,1,1,-2,1,0,0};
			139: counter1_out = '{1,0,1,1,-1,-1,-1,1,-1,0,2,-1,1,0,-1,1,0,0,2,-2,1,-1,-1,-1,1,0,2,1,-1,0,1,-1,0,0,0,-1,-1,-1,1,1,0,2,0,-1,0,0,0,1,0,0,0,-1,0,2,1,-2,2,1,0,-1,1,1,0,-1,1,0,-1,1,1,0,0,0,2,1,1,1,0,1,0,-2,1,-1,0,0,1,0,2,0,1,0,0,1,1,1,1,-1,0,0,0,-1};
			140: counter1_out = '{0,0,2,0,0,-1,0,0,0,0,0,2,-1,0,1,1,-1,0,-1,0,0,-1,2,-1,-2,-1,0,2,0,0,0,0,-1,0,-1,-1,1,-2,1,-2,-1,1,0,0,0,2,1,0,-1,-1,-1,0,0,0,-2,-1,1,2,-1,1,1,-1,0,0,-1,0,-2,0,-1,-1,0,1,-2,-1,1,1,-1,2,0,0,0,-2,-1,-1,1,1,1,0,0,0,1,0,0,0,-1,1,1,0,0,-1};
			141: counter1_out = '{0,0,1,1,1,0,0,-1,0,0,0,-2,1,0,0,-1,1,0,2,-1,-1,0,-1,0,-1,-2,1,0,-2,0,2,1,-1,0,-1,-1,1,0,0,0,-1,1,-2,1,2,-1,1,0,0,1,1,-2,1,-1,0,1,1,0,0,-1,0,1,1,1,1,1,2,0,0,0,-2,1,0,0,-1,-1,2,0,0,1,1,1,0,-1,0,1,1,1,1,0,0,0,-1,0,-2,-1,1,1,0,0};
			142: counter1_out = '{0,2,-1,-1,-1,2,0,1,0,0,0,1,0,1,0,-1,1,1,1,1,0,-2,1,-2,0,-1,0,0,0,0,-1,0,1,-1,-1,-1,3,0,2,0,1,-1,-1,0,-1,1,1,1,0,1,0,0,-1,1,-1,0,1,0,2,-1,0,0,0,-1,1,-1,1,1,1,0,-1,1,1,0,1,1,2,1,-1,2,0,0,0,-1,0,0,0,0,1,0,-1,0,1,0,0,0,0,1,-1,0};
			143: counter1_out = '{0,2,-1,0,0,0,0,1,-1,1,2,1,0,-1,0,-2,0,0,1,-3,1,1,0,0,0,-2,0,1,-1,0,2,0,0,-2,-1,-1,0,0,-1,0,0,1,2,1,0,1,0,-1,-1,1,1,0,-1,0,0,1,0,-1,-2,1,-2,-1,0,1,-1,-2,0,0,0,1,0,0,0,0,-1,1,-1,1,0,1,1,1,1,0,-2,1,1,-1,1,0,-1,1,-1,-1,0,-1,0,0,0,-2};
			144: counter1_out = '{0,0,0,1,1,-1,1,1,-2,0,-1,1,0,-1,-1,0,-1,1,-1,0,-1,0,-1,-1,-1,0,1,1,-1,2,0,1,1,0,0,-1,1,0,0,0,0,3,0,0,-1,0,0,0,0,-2,0,0,1,-1,-1,1,-1,0,-1,1,1,1,1,0,2,2,0,-1,0,0,1,1,-1,0,1,1,-3,1,1,-1,1,-1,0,1,0,1,0,-1,0,1,0,1,0,1,2,0,1,-1,0,0};
			145: counter1_out = '{-1,0,-1,0,-1,-1,1,0,0,0,-1,-1,0,1,1,0,1,0,-1,-2,-1,-1,2,1,0,0,0,1,0,1,-2,1,-2,1,1,1,-1,2,0,0,0,0,0,0,0,-2,0,1,-1,2,0,0,-1,0,0,-1,1,0,1,1,1,1,2,0,0,1,-2,0,-1,-2,-1,-1,-1,0,1,0,3,1,-1,0,0,1,0,0,1,1,0,-1,1,1,2,0,-3,1,-1,-1,1,0,0,-1};
			146: counter1_out = '{0,0,-1,-1,-1,-1,0,2,1,2,0,1,0,0,-1,-1,-1,0,-1,-1,0,1,-2,0,-1,-1,-2,0,-1,1,1,0,-1,-2,2,2,0,-1,0,-1,0,1,-1,-3,1,1,0,0,-1,1,2,-1,1,0,-2,-1,2,-2,-2,1,0,0,-1,-2,1,0,0,0,0,0,1,1,-1,-2,-1,-1,1,2,-1,1,0,1,-1,-1,0,-1,0,0,0,2,-1,0,0,2,0,0,0,0,2,1};
			147: counter1_out = '{1,0,-1,0,0,1,0,-1,0,0,2,1,-1,0,1,0,-2,-1,0,0,-2,1,1,-2,-1,-1,0,-1,-1,1,0,1,1,1,1,1,1,-1,1,1,-1,1,0,1,1,0,0,-1,1,1,-1,0,0,1,-1,0,0,2,-1,2,1,0,-2,1,2,-1,0,-1,0,0,0,1,-1,-1,1,-1,1,0,0,1,-1,2,-1,0,-1,0,0,1,1,1,0,2,-1,0,0,1,0,-1,-1,0};
			148: counter1_out = '{0,-1,0,-1,-1,1,0,2,1,1,0,1,1,0,0,0,-1,-1,2,3,0,2,2,1,0,-1,-1,0,2,0,0,0,-1,1,0,-1,0,1,2,-1,0,-1,0,0,1,-1,0,0,1,-1,0,0,2,0,0,0,-1,-1,0,0,-2,0,0,0,1,0,-2,0,0,1,0,-1,-1,0,0,-1,1,0,0,0,0,-2,1,1,0,0,-1,0,0,0,1,-1,1,0,0,-1,0,-1,0,0};
			149: counter1_out = '{-2,0,-1,0,0,0,0,0,0,-1,-1,1,0,0,0,1,0,0,0,1,1,2,-1,0,-1,0,0,3,2,1,1,-1,-1,0,0,-1,-1,0,0,0,-1,-1,-1,-1,2,0,1,0,-2,-1,-1,-2,-1,0,0,-1,0,0,-1,0,2,1,-1,-1,0,0,1,-1,0,0,1,0,1,0,2,0,1,-2,1,-1,0,0,2,1,0,0,1,-3,0,-1,-1,1,2,0,-1,2,0,-1,0,1};
			150: counter1_out = '{1,-3,0,-1,0,-1,-1,0,1,0,1,1,1,0,2,0,-2,-1,-1,-2,1,1,0,2,1,1,1,-1,1,1,2,-2,1,0,1,-1,-1,-1,2,2,-1,-2,0,0,2,-1,-1,0,1,0,0,-1,0,0,2,0,2,-1,0,0,0,0,-1,2,2,-1,0,0,1,1,-1,0,-3,-1,1,0,2,0,-1,-2,0,0,1,-2,1,-1,0,-1,-1,-1,-1,0,-1,-1,-1,0,0,1,0,-1};
			151: counter1_out = '{-1,-2,-1,0,0,-1,-1,1,-2,1,1,1,1,-1,-1,1,1,-1,0,-1,-1,2,0,-1,-1,0,0,2,-1,-1,1,1,2,-1,0,1,-1,-2,0,0,-1,0,0,0,0,-1,0,0,-2,0,-1,-1,-1,-2,-1,-1,0,2,0,-2,-1,-1,0,-2,1,1,0,-1,1,-1,-2,1,0,0,0,0,1,0,1,0,0,1,1,-1,3,0,-4,-3,-1,0,1,0,1,0,-2,1,0,-1,0,-3};
			152: counter1_out = '{1,0,0,0,-1,0,2,-1,0,0,-1,1,1,-1,-1,0,1,0,1,-1,-1,0,0,1,-1,-2,0,1,1,0,3,-2,2,0,0,2,-1,-2,0,0,0,0,-1,-1,0,-1,1,-1,0,1,-1,-1,0,-1,-1,-1,1,0,1,-1,-1,1,3,0,0,0,-2,-1,1,0,-2,0,0,-1,0,2,1,1,-1,-1,-1,0,0,1,2,-1,-1,1,0,0,-1,0,-1,0,-2,0,2,0,-1,1};
			153: counter1_out = '{-1,1,0,-1,0,0,0,1,-2,-1,-1,1,1,-2,0,1,1,-3,0,-1,0,0,0,0,1,-1,0,2,-1,0,-1,-1,2,1,1,1,-1,1,0,0,0,0,0,2,0,1,-1,0,0,-1,1,-2,2,0,-1,-1,-2,1,-1,1,-2,1,0,-1,0,1,-2,-1,0,-1,-1,0,3,-1,0,1,0,1,1,0,-3,0,0,-1,1,-1,-1,-1,-1,-2,-2,-1,-1,-1,-1,1,0,-1,0,1};
			154: counter1_out = '{1,-1,-2,0,-1,-1,0,1,0,2,-2,2,0,0,-1,0,0,-2,0,1,-2,1,0,1,1,0,0,1,-1,-1,1,0,0,1,0,0,-3,-1,-1,0,0,-1,0,1,0,1,-1,1,1,-1,-1,1,0,1,1,-3,1,-2,-2,-1,-2,0,-2,0,1,-1,1,1,0,0,-1,1,1,1,0,-1,0,-1,1,0,1,0,0,1,0,1,-1,-1,0,0,0,1,-1,1,-2,0,2,1,0,2};
			155: counter1_out = '{-1,1,-1,-1,0,-1,2,1,-1,0,-1,-1,1,-2,-1,2,0,-1,-1,-1,0,1,-2,0,-1,0,0,2,-1,1,0,-1,-1,0,1,1,0,1,-1,1,0,0,-1,0,1,0,1,0,0,0,0,0,2,0,0,-1,-1,-2,-1,0,1,-1,-1,-2,-1,-1,0,1,0,-2,-1,0,1,-2,1,-2,0,0,1,2,-1,1,0,-2,-1,-1,0,1,0,-2,0,-1,-2,0,-1,0,1,1,-1,1};
			156: counter1_out = '{1,0,0,-1,-1,-2,1,0,1,1,-2,0,-1,0,0,0,0,0,-2,0,-1,0,1,1,0,-1,-1,-1,0,-1,1,-1,0,0,2,2,-2,-1,1,1,0,0,0,0,1,0,-1,-1,-1,0,-2,0,1,0,1,0,-1,1,-1,1,-1,0,-1,1,-1,1,0,0,1,0,-2,-1,0,-2,1,2,2,1,2,-1,0,-1,0,0,-1,0,0,0,0,0,0,0,-1,-2,-2,1,1,0,0,0};
			157: counter1_out = '{-1,1,-2,1,0,1,-2,1,0,0,-1,1,0,1,0,0,1,-1,-2,-1,-2,-1,-1,0,-1,1,1,1,0,0,0,0,0,-1,0,0,1,0,-2,0,0,1,-2,-2,1,-1,1,-1,0,0,0,0,0,-2,0,1,0,-1,0,0,0,2,1,0,0,2,0,-1,-1,1,-1,-1,0,-1,-1,-3,1,1,-2,2,-1,0,0,2,0,-1,0,1,1,0,0,-2,-1,1,-2,1,0,1,0,4};
			158: counter1_out = '{2,-1,-1,0,1,0,1,-1,0,-1,-2,1,1,0,1,0,0,1,0,0,-2,0,0,-3,-1,0,0,2,-1,1,0,-2,0,0,0,0,1,0,0,1,3,-1,0,0,0,-2,-1,-1,-3,-1,-2,1,1,-1,0,0,0,2,0,1,1,0,0,2,1,-1,1,-1,2,1,-2,0,-2,0,0,0,1,0,-1,2,1,0,1,0,0,-1,0,0,0,1,1,-1,0,1,-2,1,0,-1,0,1};
			159: counter1_out = '{1,0,-1,0,0,0,0,2,0,-1,0,1,1,2,0,1,2,1,1,1,-1,-1,2,0,-1,1,0,2,0,-1,0,-1,0,-2,-1,1,0,0,1,1,1,2,-1,0,0,-3,-1,0,0,-1,3,1,0,-1,-1,1,1,0,-1,0,0,-2,-1,1,1,0,0,1,0,-1,0,-1,-1,-1,1,0,0,-1,0,1,0,1,1,1,0,-1,-1,0,0,-1,-1,0,0,0,-1,1,0,2,1,0};
			160: counter1_out = '{0,1,-1,-1,0,1,0,0,0,-1,2,0,1,-1,0,-1,0,0,1,-1,-1,-2,0,0,1,-1,0,0,0,0,0,2,-1,1,1,1,0,1,-1,-1,-2,1,2,-2,2,0,-1,0,-2,1,0,0,1,0,1,2,0,0,1,-1,-3,-1,-1,-1,0,1,3,0,-1,0,0,1,-2,0,0,1,-1,0,0,1,-1,1,-1,0,0,0,0,0,-1,0,1,-1,-1,1,-1,0,1,1,1,0};
			161: counter1_out = '{-1,0,0,0,-1,-2,2,-2,-1,-1,2,1,1,0,0,-2,2,0,0,-1,0,-1,1,1,-1,0,1,0,0,0,-1,-1,-1,1,-1,-1,-2,-1,0,1,-2,1,0,1,0,0,0,0,-1,-1,-1,-2,1,2,-1,-1,-1,1,-1,0,1,1,-1,1,-1,1,1,0,1,-1,1,1,0,0,0,0,0,0,0,2,0,0,1,-1,0,-1,0,1,-1,0,0,-2,-1,-1,1,1,0,-1,2,-2};
			162: counter1_out = '{1,-1,0,-1,-2,0,1,-2,0,2,1,1,0,1,-1,0,-1,-1,-1,-1,0,1,-1,0,-2,1,-1,0,0,0,2,0,0,0,0,-1,1,0,-1,-1,-1,1,0,0,0,0,0,0,-1,-1,1,2,-1,1,1,1,-2,0,-1,-2,-1,0,1,-1,0,1,-1,0,-1,1,1,1,0,-1,-1,0,0,1,1,-1,1,0,1,-1,1,0,1,0,2,2,0,-3,2,0,0,1,-1,1,1,-2};
			163: counter1_out = '{0,2,-1,1,-1,-1,0,-1,1,-1,-2,0,0,0,-1,0,1,2,-2,-1,0,-1,-1,1,0,1,0,-1,1,1,2,0,0,0,-2,1,2,2,-2,1,1,1,0,-1,-2,1,-2,-1,-1,1,2,1,0,-1,0,1,0,-1,-1,0,0,1,1,1,0,-1,0,0,1,-1,0,1,1,-2,1,1,1,0,0,1,0,-1,0,0,-1,0,1,1,0,1,-1,0,1,-1,-1,2,0,-1,1,-2};
			164: counter1_out = '{0,1,0,0,1,-1,1,0,-1,-1,0,0,-1,1,1,2,1,1,0,1,0,-1,-1,1,-1,3,-2,0,1,-1,0,-1,0,1,0,-2,0,0,-1,3,-1,1,0,0,-1,0,0,0,2,1,1,2,2,2,-2,1,1,-2,0,0,0,1,0,0,-1,0,0,1,0,1,1,-2,0,-1,0,1,0,0,1,-1,0,0,1,1,2,-1,-1,1,1,1,0,3,2,1,2,0,-1,0,1,-3};
			165: counter1_out = '{3,0,1,1,0,1,0,1,0,-2,-1,2,1,-1,-2,0,0,1,1,-1,-1,1,1,2,-1,-1,1,0,1,0,0,0,1,1,0,1,1,0,-1,-1,1,-1,-1,-1,1,-1,-1,0,0,-1,1,-1,-1,-1,0,1,0,-1,0,1,-1,0,0,0,0,1,-1,0,-2,-1,-1,0,0,0,-2,1,-1,1,1,0,0,2,-2,-2,0,-1,-1,0,0,1,1,1,-1,1,-1,-2,-2,0,0,-1};
			166: counter1_out = '{0,1,1,0,1,0,-1,0,1,2,1,-1,2,0,-1,0,-1,-1,1,-1,1,-1,-1,-2,0,0,-1,-1,0,1,1,-2,-1,0,-1,2,0,-1,0,0,-1,0,0,0,0,1,2,0,0,-1,-1,0,0,1,0,0,0,-1,0,-1,-1,0,1,0,1,0,1,0,0,1,-1,1,1,0,-1,-1,0,1,-1,-1,-1,-1,-2,0,0,1,0,3,0,0,1,-3,0,2,-1,-1,-2,-1,0,0};
			167: counter1_out = '{1,-1,0,1,0,0,1,1,0,1,-2,1,-2,1,2,1,0,-1,0,-1,-1,0,0,-1,0,0,1,1,1,-2,-1,1,-1,3,1,1,0,2,2,0,1,1,0,-1,0,0,-2,0,-1,3,0,-1,0,2,0,0,0,1,-2,-1,0,0,0,0,-1,1,0,-1,1,0,1,0,0,0,-1,1,0,0,0,1,1,1,-1,2,0,-1,-1,0,-1,-2,-2,1,1,-1,0,0,-1,1,1,0};
			168: counter1_out = '{0,0,-1,1,1,0,0,-1,-1,0,2,-2,1,2,0,2,-1,-2,-2,-1,-1,0,-1,0,-1,1,1,-1,-1,0,-1,1,-1,-2,0,2,0,0,0,0,2,0,0,0,2,0,1,1,-1,-1,0,1,-1,0,0,1,0,-1,0,-1,1,0,0,1,-1,1,-1,-1,1,1,0,0,-1,2,0,-1,-2,0,0,1,-1,1,-1,0,1,1,1,2,-1,1,0,-1,-1,0,0,-1,0,0,0,-2};
			169: counter1_out = '{-1,0,0,0,0,-2,1,0,0,1,-2,-1,-2,0,1,1,0,-1,1,0,0,0,-1,0,-1,0,0,0,2,0,0,0,1,-1,0,1,-1,2,0,-1,1,0,0,-1,-1,-1,-1,-2,1,-3,-1,0,1,-1,0,-1,2,0,1,0,0,-1,0,0,-1,1,0,0,-1,-1,1,1,-1,-1,1,0,-1,1,1,-1,-1,-1,-2,0,0,1,1,0,-1,-1,-1,2,1,2,-1,0,1,0,0,0};
			170: counter1_out = '{0,1,1,-1,2,-1,1,2,2,0,0,0,-1,2,1,0,1,1,0,1,-1,-1,1,0,1,0,0,-1,0,-1,2,0,1,1,-3,-1,1,-3,1,2,-1,1,-1,2,-2,0,0,-1,0,0,1,0,-1,-1,0,1,0,0,-1,-1,0,0,0,-1,0,0,1,0,-1,2,0,-1,1,0,0,1,-1,0,1,-1,1,2,0,0,1,0,-2,0,-1,0,1,0,0,0,1,0,3,-1,0,0};
			171: counter1_out = '{1,-1,-2,0,-1,1,-2,-1,2,-1,2,3,0,1,2,1,-1,-1,0,-1,0,0,1,1,-1,-1,2,-3,1,0,-2,-1,0,0,0,0,-1,0,-2,1,0,-1,1,-2,0,0,1,-1,-1,-1,-1,1,1,1,-1,1,0,1,1,1,-1,1,2,1,0,0,1,-1,1,1,-1,0,0,0,0,1,0,0,0,1,-1,1,-1,1,1,1,-1,1,-1,0,1,-1,-1,0,0,0,-1,-2,1,-1};
			172: counter1_out = '{0,-1,0,-1,-1,0,0,0,-1,0,1,-1,0,0,1,1,2,-1,1,0,3,-1,-1,0,1,-1,0,0,1,0,0,-2,0,1,1,2,0,3,2,0,-1,1,-1,1,-1,0,-1,0,0,1,0,0,0,0,-1,0,2,-1,0,0,1,0,-1,-1,0,-1,-2,0,-1,0,-2,1,0,0,0,0,-1,0,1,1,0,1,0,2,0,0,1,1,0,0,0,0,1,-1,-1,-1,0,1,-1,0};
			173: counter1_out = '{0,-1,2,0,-1,1,-2,0,0,-1,1,-1,0,1,-1,2,0,0,-1,0,0,1,1,2,0,1,2,3,-1,1,2,-1,1,-1,-1,-1,3,0,1,-1,-1,-1,2,1,0,-1,-1,1,2,0,1,0,0,0,2,1,0,1,0,0,-1,2,-1,0,1,2,0,2,1,2,-2,-1,-1,0,2,-1,1,-2,-1,-1,0,0,0,1,1,0,-1,-1,0,1,-1,0,0,-2,0,0,0,1,0,0};
			174: counter1_out = '{1,1,1,-1,1,0,-2,1,1,0,3,2,0,1,0,1,-1,0,-2,1,1,1,1,-1,2,-1,0,-1,-1,0,0,-1,0,-1,2,0,0,1,1,1,-1,2,-2,2,0,0,0,2,0,1,2,-1,0,2,-2,1,1,0,0,0,0,0,2,0,-1,0,1,-2,0,-1,0,1,0,0,1,0,1,-2,-1,0,1,1,0,1,-1,-2,2,0,2,1,0,1,0,-1,0,-1,-1,0,-2,-4};
			175: counter1_out = '{0,1,-1,1,-2,0,1,1,-1,0,0,-1,2,1,-2,1,0,0,0,1,0,1,0,1,-1,0,0,-1,2,0,0,-1,0,2,-1,0,-1,-1,2,0,1,1,1,0,1,-1,0,0,-2,1,1,-2,0,-1,-1,-1,-1,0,0,0,0,0,1,-1,-1,-1,-2,0,1,-2,0,0,-2,0,0,-1,-1,1,0,-1,1,0,1,-2,-1,-1,1,0,1,-1,2,-2,0,-2,-1,1,-1,0,1,-1};
			176: counter1_out = '{1,0,1,-1,0,0,-1,0,0,1,-1,-1,1,0,0,1,0,1,0,0,-1,0,1,2,0,0,-1,2,0,-1,0,-1,1,0,0,-1,1,-1,2,0,1,0,1,-1,1,0,0,0,0,0,1,1,-1,-1,-1,-1,2,1,-1,-1,2,-1,1,0,0,0,-1,1,2,1,-2,1,0,0,2,0,0,-1,0,-2,-1,0,1,-1,-1,2,0,0,-2,-1,0,0,2,-1,-2,0,1,1,-2,0};
			177: counter1_out = '{1,1,1,1,0,1,0,1,-2,2,-1,0,0,-1,0,0,-1,1,-1,-2,0,1,-1,0,0,0,0,2,0,-2,-2,0,1,0,2,1,0,-2,3,1,1,0,-3,1,0,-2,-1,1,2,-1,1,0,0,1,-2,0,2,0,-1,1,0,1,-1,1,1,2,1,-1,1,1,-1,0,1,0,0,-1,2,-3,3,-1,1,-1,0,-1,-2,0,3,-1,0,0,1,-1,0,-2,-1,1,-1,1,0,-2};
			178: counter1_out = '{-1,0,0,0,-2,0,0,-1,2,0,-1,1,-1,1,0,-1,-2,1,1,-2,0,1,1,0,0,-1,-1,1,0,0,-1,0,0,0,1,-1,-1,0,0,-1,1,-2,-1,-1,0,1,-1,2,0,2,2,0,0,-3,0,-1,2,-1,0,1,-1,-1,2,-1,1,1,1,0,2,0,0,-3,-1,-1,1,0,0,-2,1,0,2,-1,1,0,0,1,1,-1,-2,0,-1,-1,1,0,-2,1,0,2,0,1};
			179: counter1_out = '{2,-2,-2,-1,-1,-1,0,-1,-1,2,1,1,0,-1,0,1,-1,0,0,-2,-1,-1,2,1,-2,0,-1,0,-1,0,-2,2,1,-1,-1,0,1,0,0,0,0,0,1,0,0,1,0,1,2,-1,-2,1,-2,0,-1,-1,-1,-1,-1,0,0,-3,0,0,0,-3,0,1,2,0,0,0,-1,1,0,2,1,0,1,-1,1,-1,0,-1,-2,0,1,-2,0,-2,0,1,1,0,1,0,0,-1,1,0};
			180: counter1_out = '{-1,0,-2,-2,1,0,2,0,0,0,-1,0,1,-1,0,0,0,-2,-3,-1,0,0,0,-1,-1,0,0,0,-1,0,2,2,-1,-1,-1,-2,-2,0,1,0,0,1,-1,-1,0,0,1,1,0,0,0,0,-1,-1,0,-1,0,-1,0,1,0,-2,0,-1,1,3,3,1,1,1,-2,-3,-1,1,-1,-1,0,-1,0,-1,0,0,0,0,-1,-1,0,0,0,-1,-1,0,-1,1,1,-1,0,-1,1,-1};
			181: counter1_out = '{1,1,0,0,-1,0,2,1,0,0,-1,0,1,-1,-1,1,1,-2,-1,-1,0,-1,0,-1,1,0,0,2,0,0,0,1,0,1,1,0,0,-1,0,1,1,0,-1,0,0,0,0,-1,0,0,1,0,0,0,0,-2,-1,1,-1,1,1,-1,-1,-2,1,-1,-1,-1,-2,2,-2,1,-2,-1,0,0,2,0,1,-2,0,2,1,-2,0,0,-1,-3,-1,-2,1,-1,-3,-1,0,-1,1,-1,1,0};
			182: counter1_out = '{1,-1,0,1,1,3,1,0,0,-1,1,2,1,-1,-1,1,-1,-3,1,-1,-1,0,0,-1,-2,1,0,1,1,-1,-1,1,2,1,0,1,-1,0,-1,0,0,0,0,-1,0,0,0,-1,0,1,2,0,0,1,0,-2,1,0,0,-2,-1,1,-2,0,1,-1,0,0,0,0,-2,0,0,0,1,1,0,1,0,0,0,2,-1,2,1,1,0,0,2,-2,0,-1,-1,0,0,3,1,-1,-1,0};
			183: counter1_out = '{0,0,3,0,0,1,2,1,0,0,-1,-1,-1,0,1,1,0,-1,0,-1,-1,-1,1,0,1,-1,1,0,0,1,0,-1,0,2,-1,0,-1,-1,0,-1,1,-2,0,1,1,0,-1,1,0,0,-1,2,-1,-2,0,0,1,-1,-1,-2,0,-1,-1,1,0,1,0,0,2,1,-1,0,1,0,-2,-1,0,0,0,-2,0,2,1,-1,0,-1,-1,1,0,-1,1,-1,-1,0,0,1,2,1,1,1};
			184: counter1_out = '{1,0,1,1,-2,4,-2,1,-1,1,0,0,0,0,-1,0,0,-1,1,0,1,1,0,-1,-1,1,1,1,0,0,-1,0,0,1,-2,0,-1,-2,0,-2,-1,1,-1,-1,0,-1,-1,0,0,-1,1,-1,-1,0,0,-1,0,0,-3,0,2,-1,1,0,-1,0,0,-1,0,0,-1,0,1,0,1,0,1,0,0,1,0,0,-1,0,0,-2,1,0,-3,-1,-1,0,-1,-1,-1,-1,1,0,-1,2};
			185: counter1_out = '{0,-1,-1,-1,-1,0,-2,-1,-2,1,2,0,0,1,0,-1,1,0,0,0,1,2,2,-2,1,1,2,-1,-1,0,1,-1,1,0,-2,0,1,-1,-1,-1,-1,1,0,2,1,0,-2,1,1,1,0,0,0,-1,0,-2,0,2,-2,0,0,0,-1,0,-2,-2,2,-1,1,-1,1,1,1,1,-1,0,-1,1,1,1,0,5,-1,-1,-1,1,0,0,-1,0,1,1,0,-1,0,-1,1,1,0,3};
			186: counter1_out = '{1,0,0,0,1,1,-2,0,-1,-1,2,1,0,0,0,1,1,2,0,0,0,-2,0,-1,-1,-1,1,0,0,0,0,-1,1,0,-1,-1,0,-1,0,0,1,0,-1,-1,1,2,-1,-3,-1,-1,2,0,1,0,0,1,1,-1,1,0,-1,-1,-2,0,0,1,2,-1,1,-1,0,0,-3,1,-1,-2,0,-1,0,0,1,1,0,0,0,-2,0,0,-2,1,1,-1,-2,-1,1,-1,0,0,0,1};
			187: counter1_out = '{0,1,0,0,-1,1,-2,-1,-1,1,1,0,1,-1,1,1,1,0,0,0,1,-2,1,2,1,2,1,1,-1,1,2,1,-2,1,1,0,2,0,0,0,0,0,0,0,0,-2,1,-1,-1,1,0,1,0,-1,1,0,1,0,1,-1,0,1,-1,-1,-2,0,2,-1,1,0,1,-2,-1,-1,1,1,0,2,2,1,-1,1,0,0,1,-1,0,-1,0,1,0,-1,1,-1,1,-1,1,0,2,0};
			188: counter1_out = '{0,-1,-1,1,-1,1,1,0,-2,0,2,2,-1,0,0,0,2,1,1,-1,0,0,0,0,0,0,0,2,2,-1,0,0,-2,-1,3,1,0,1,-2,-1,-1,0,0,-1,0,1,-1,0,0,-1,0,0,-1,0,0,0,0,-1,0,0,-1,0,-2,0,-1,0,3,0,1,-1,-1,0,-1,0,-1,2,0,0,1,0,0,0,-2,2,0,-2,0,0,-1,0,0,-1,-3,-2,0,0,0,1,1,-1};
			189: counter1_out = '{-2,0,-1,-1,2,0,1,1,1,0,1,-1,0,1,2,-1,0,1,-1,-1,-1,0,0,-1,0,1,-1,1,-1,0,-1,0,1,1,-1,1,-3,0,-1,0,-2,0,0,0,-2,1,1,0,0,0,0,0,1,2,1,0,2,1,-2,0,-1,-1,-1,1,0,-1,0,-2,1,-1,1,-1,0,0,0,0,-1,0,0,0,0,-1,1,0,-1,0,1,1,-1,0,0,0,0,0,0,-2,0,1,1,-2};
			190: counter1_out = '{0,-1,0,0,-1,1,2,0,0,0,1,2,0,-1,-1,-2,-2,0,0,-1,1,0,0,-2,1,0,1,2,0,1,-2,1,0,1,0,-2,0,-1,-2,-1,1,2,0,-2,0,-2,1,1,0,2,-1,-1,-1,-1,0,-1,0,0,1,-1,-1,0,0,0,1,1,1,0,1,1,-1,1,-2,0,1,0,2,1,-1,2,1,-1,0,0,0,0,-2,-1,0,0,0,2,-1,0,1,0,-1,2,0,-2};
			191: counter1_out = '{1,0,-2,0,-1,-1,1,2,-2,1,0,2,-1,0,0,0,1,-2,0,1,1,1,-1,1,-2,1,0,0,1,1,1,1,-2,-1,0,0,0,1,-2,-1,-1,2,-1,-1,0,-1,2,1,-1,-1,-1,0,-1,-1,-1,0,0,1,-2,1,-2,0,-1,-1,2,0,1,0,-1,1,1,0,-1,-3,0,0,2,1,0,-1,-1,-1,1,1,0,-1,2,-1,-1,0,-1,-1,0,0,0,1,0,2,1,-2};
			192: counter1_out = '{0,0,0,0,1,0,1,-1,1,2,0,-2,0,-2,-4,0,0,0,2,0,-1,-1,0,0,-2,-1,0,-1,1,0,0,1,-2,-1,1,-1,-2,2,-1,2,0,-1,1,0,0,0,0,-1,0,2,0,-1,-1,0,1,1,0,0,1,-2,-3,-1,-1,0,-2,-1,0,0,2,1,-1,-1,1,1,-2,-1,0,1,0,0,2,0,0,1,1,-1,1,1,-2,2,1,0,1,0,-1,-1,-1,0,1,-1};
			193: counter1_out = '{0,0,-1,1,0,2,1,0,-2,0,-2,-1,-1,0,-1,0,-1,0,-1,-2,0,1,-1,0,0,-1,0,0,0,0,1,1,-2,0,1,-1,0,0,-1,1,-1,0,2,1,1,-1,0,-1,0,1,-1,-2,1,-1,-1,1,1,1,-1,-1,1,-1,0,0,1,0,-1,0,-2,2,1,-1,1,-2,1,-1,0,0,1,0,2,-1,0,-2,0,-1,2,-1,0,1,0,-3,0,0,-1,-1,0,1,-1,1};
			194: counter1_out = '{0,0,0,0,0,-1,1,1,1,-2,0,-2,0,0,1,0,0,-1,1,0,0,-2,-1,-2,-2,0,0,1,-1,1,-1,-1,1,0,-2,-1,0,1,-2,-2,1,0,-4,0,0,1,1,0,-1,1,-1,0,-3,-1,0,0,0,1,-2,0,0,0,-1,0,0,0,0,0,-1,1,-1,0,0,-1,0,-2,2,-1,1,-1,1,1,-1,0,0,-1,-1,2,0,0,0,0,0,-1,0,0,1,0,0,1};
			195: counter1_out = '{-1,1,1,1,1,0,0,-2,0,-1,-1,-2,-1,0,0,-1,0,-1,-1,1,2,0,1,-1,1,1,2,-1,1,-1,0,0,1,1,0,-1,0,0,-1,1,-1,0,2,-1,0,-2,-1,2,-1,0,0,-2,0,1,2,0,-1,-1,1,-2,-1,0,-1,0,-1,0,-1,0,-1,-1,-2,0,-2,1,-1,1,-1,0,-2,-1,0,-1,1,0,1,0,-1,0,1,-1,0,-1,1,2,-1,0,0,-1,0,1};
			196: counter1_out = '{-3,0,-1,2,-1,1,0,-1,-1,0,-1,-1,2,-1,-1,-1,-1,0,-2,2,0,0,-1,0,-1,0,-2,1,-1,-1,0,-2,1,1,1,-1,-1,-1,-1,-1,2,-1,-1,0,0,1,0,1,-1,-2,-4,-3,3,1,3,0,-1,-2,1,0,0,1,1,0,1,0,0,1,0,0,0,-1,-1,-1,0,0,0,-1,1,1,2,-1,-2,0,1,1,2,-2,1,0,1,1,0,1,-1,-1,0,1,1,1};
			197: counter1_out = '{1,0,0,0,-1,0,2,-1,0,-2,1,2,0,-1,-1,-2,3,0,-1,1,1,1,-2,0,1,0,1,0,0,-2,-1,1,-1,-1,-1,2,1,1,1,0,0,0,0,0,0,0,0,1,3,-1,0,1,0,2,0,0,0,1,1,2,1,2,0,0,0,-1,0,1,0,0,0,-2,0,0,2,0,0,-1,0,2,1,0,0,2,0,2,0,2,-1,-1,-1,1,0,1,0,0,-1,-2,1,-1};
			198: counter1_out = '{0,2,1,0,1,1,-1,0,0,0,-3,1,-1,0,0,0,2,1,0,-1,-1,0,1,1,0,3,0,-2,2,0,2,2,1,0,0,0,0,0,1,0,1,1,1,1,-1,1,0,0,1,-2,1,1,-1,1,-1,1,0,0,0,-1,0,1,-1,-1,0,-1,0,0,0,0,0,0,1,1,-1,0,0,0,0,0,2,-2,1,-1,0,-1,2,0,0,-1,1,0,1,0,0,1,0,-2,-1,-1};
			199: counter1_out = '{1,0,0,1,0,1,0,-1,1,0,1,-1,0,1,-1,0,1,0,-1,0,1,0,-2,0,1,-2,-2,0,0,1,0,-1,-1,0,1,-1,0,2,-3,-1,1,0,0,-1,1,0,0,2,2,-1,-1,-1,-1,0,0,1,1,1,1,-1,0,1,0,0,0,1,0,0,0,-1,0,1,-2,0,3,-1,0,1,-1,0,1,0,0,1,-1,0,2,2,1,0,-1,0,0,1,-1,1,0,-1,-1,1};
			200: counter1_out = '{0,-1,-1,0,0,0,-2,-1,-1,-1,-1,1,1,-1,1,-1,1,-2,0,1,0,1,-1,-1,1,0,1,-1,-1,0,0,-2,-1,1,1,-1,0,0,1,1,0,0,1,-1,-1,0,2,-2,0,-1,-1,-1,0,0,0,1,0,1,1,-1,-1,-3,-1,0,0,0,-2,0,0,1,0,1,0,1,0,-1,-1,1,0,1,0,1,-1,-1,0,1,-2,-1,-1,0,-2,0,2,0,0,1,0,1,1,-2};
			201: counter1_out = '{1,1,1,-1,2,1,-1,1,1,0,1,-1,0,-1,0,0,-2,0,0,2,-1,2,1,0,1,-1,0,0,1,2,1,1,1,1,0,0,0,2,-1,1,0,0,0,1,1,3,-2,-1,1,2,0,2,-1,0,1,1,-2,1,0,-1,1,0,-1,2,0,-1,-1,2,0,-1,0,-1,0,1,1,-2,0,1,-1,1,-1,0,-1,2,0,-1,1,-1,-3,1,-1,0,1,1,-1,1,1,-1,-2,-1};
			202: counter1_out = '{1,1,0,0,2,0,-1,-1,0,1,-1,1,0,-1,-1,2,1,2,0,1,1,2,0,2,1,-1,0,-1,0,0,1,0,1,1,2,-1,-1,-1,3,0,-1,1,-1,0,2,0,-1,0,1,1,1,-1,0,1,-1,-2,-1,1,-1,-1,1,1,0,-1,1,-2,-1,0,0,1,2,1,-1,-1,-1,1,0,0,0,2,-1,-1,0,0,2,-1,-1,-2,-2,1,1,-1,1,2,-1,0,1,0,0,0};
			203: counter1_out = '{0,1,-1,0,0,1,-1,2,-1,0,0,-1,-2,-1,1,1,-1,1,-2,2,0,0,-1,3,1,-1,0,-1,1,0,-1,-1,2,0,0,0,-1,1,1,0,0,0,-1,1,1,-1,-1,-1,0,2,1,1,0,1,-1,-1,-2,0,-1,-1,-1,0,1,0,0,2,-1,-2,0,-1,1,0,-1,1,-1,0,0,0,-1,0,-1,-2,0,1,1,-1,0,0,0,-1,1,-1,-1,1,1,1,0,0,0,0};
			204: counter1_out = '{1,-1,0,0,0,-1,0,-1,-1,0,-1,1,1,1,0,0,0,2,0,0,1,3,1,-1,-1,-1,1,0,0,0,0,-1,0,2,-1,-1,2,0,3,1,-2,2,1,1,0,0,1,1,-1,-1,0,-1,1,0,-2,1,1,1,-1,1,0,-2,-1,0,1,0,1,0,1,1,0,-1,-1,1,-1,-1,0,0,1,1,1,0,1,-2,0,-2,1,-1,1,-3,0,1,1,0,0,1,1,2,-1,0};
			205: counter1_out = '{1,-2,1,0,-1,0,1,0,0,2,0,0,-1,-2,0,0,0,0,0,0,0,0,1,-1,1,1,0,0,0,-2,0,-1,1,1,0,-1,0,-1,1,0,1,-1,1,0,1,0,1,0,0,0,-1,-1,1,-1,-1,0,1,1,0,0,-1,0,0,-1,1,-1,1,-2,-1,-2,2,-3,0,1,-1,0,0,-1,3,1,0,-1,1,0,-1,-2,2,1,0,1,-1,0,2,0,1,2,0,-1,1,-1};
			206: counter1_out = '{1,-1,-1,-1,-2,0,-1,0,0,1,1,1,1,0,0,1,0,0,-1,0,0,1,-1,0,0,0,0,0,1,0,-2,1,0,-1,0,-1,0,-1,0,0,-1,1,-2,0,-1,1,-1,-1,0,-1,1,-1,-1,-1,0,-1,0,0,-1,0,0,1,0,0,1,2,0,-1,2,0,2,0,-3,1,0,0,2,0,1,1,-1,-1,1,1,1,0,2,0,-1,1,-1,0,1,0,0,2,0,0,-2,-1};
			207: counter1_out = '{0,-1,-1,-1,1,1,1,-1,0,1,-1,0,-1,0,1,0,0,0,1,0,-1,0,1,-1,0,-1,2,0,2,1,-1,-1,1,0,-1,-1,0,0,-2,0,-1,1,-2,1,-1,0,0,2,0,1,0,0,-1,0,-1,-2,0,1,-1,2,0,-1,1,-2,1,1,-1,0,3,-1,1,0,1,0,-1,1,0,-1,1,-1,0,-3,3,-1,-1,1,0,0,0,-1,1,1,1,0,0,-1,1,1,0,-1};
			208: counter1_out = '{2,-1,0,0,1,1,0,0,1,2,-2,1,0,-1,1,0,0,0,0,-2,-1,-1,1,-2,1,0,0,-1,0,1,-1,0,-3,2,0,1,0,0,-1,0,0,0,-1,2,0,2,-1,-1,1,0,1,0,-1,-1,1,-1,2,1,0,-1,0,0,1,-1,1,1,0,-2,0,0,0,-1,-1,-1,0,0,0,1,1,0,1,-4,0,0,0,-1,0,0,-2,-3,0,-1,0,0,0,0,2,3,0,0};
			209: counter1_out = '{0,-1,-1,-1,1,1,0,0,0,0,-1,1,0,1,-1,2,-1,-3,0,-3,0,1,2,0,0,-1,0,-2,-1,2,-2,1,0,0,-1,1,-1,0,0,0,-1,-1,-2,-2,0,0,0,-2,-1,1,-2,-1,2,0,-2,-1,0,1,0,1,-1,-2,1,1,0,0,-2,1,0,1,1,0,-2,0,1,-1,1,-1,-1,-2,0,-1,0,0,-1,-1,1,0,-1,0,-1,1,1,-1,1,0,0,4,1,-2};
			210: counter1_out = '{2,2,-1,1,0,1,1,0,1,1,0,-1,-1,0,-1,1,-1,-3,-2,-1,0,0,1,-1,-1,0,-1,-2,1,-1,0,-1,-1,0,0,0,-2,-1,-1,1,1,-3,0,1,0,0,0,-1,-1,1,1,-2,1,-1,2,-2,-1,0,0,1,0,0,-1,-1,-2,0,0,2,0,2,1,-1,1,-1,1,0,-1,0,0,-2,1,-1,2,0,1,0,-1,1,0,-1,0,-1,2,-1,-2,0,0,2,0,1};
			211: counter1_out = '{0,-1,1,0,1,3,0,1,-1,0,3,2,0,0,-1,-1,2,-1,-2,-1,-1,-1,1,0,-2,-1,-1,1,-2,-1,1,0,-1,2,1,0,-1,-1,-1,2,0,-1,0,-1,0,2,0,-1,-1,-1,1,1,-1,-1,-2,-2,1,0,0,-3,0,0,-1,-1,-1,1,-1,-1,0,2,0,-1,2,-1,1,0,1,0,-1,0,-1,3,-1,0,-2,0,1,0,2,0,1,2,1,-2,0,0,0,1,-1,1};
			212: counter1_out = '{0,-1,1,1,-1,1,1,0,1,-1,0,2,2,1,0,0,0,1,0,-2,0,1,0,0,0,0,-1,2,0,-1,0,-1,-2,1,-1,1,1,-1,0,0,0,0,0,-1,-1,1,1,-2,-1,1,2,0,1,1,1,-1,1,1,0,-2,0,-1,-1,-1,-1,2,-1,1,-1,0,1,3,0,0,-1,-2,1,2,3,0,0,1,2,-1,-3,0,0,0,0,-1,-1,1,0,0,0,-2,0,2,0,2};
			213: counter1_out = '{1,1,0,0,0,3,-2,0,0,0,1,1,2,0,0,0,1,2,0,0,0,0,0,0,0,0,1,0,1,2,2,-1,0,-1,-1,0,1,1,1,-1,0,-2,-1,1,-1,3,1,-3,0,0,1,1,1,-1,0,1,0,-2,0,-1,-2,-1,0,2,0,-1,1,0,2,1,0,-1,0,1,-1,1,1,-1,-1,2,-1,-2,-1,0,0,1,0,0,-1,0,0,-2,-1,0,-1,0,1,0,0,4};
			214: counter1_out = '{1,-1,0,0,0,1,-3,0,1,1,2,1,0,0,0,0,1,0,1,-1,0,2,-1,1,0,2,1,2,0,2,0,0,-2,-1,1,0,1,1,0,1,-2,0,1,0,0,2,-1,-2,1,0,0,0,1,0,1,0,1,0,1,-1,0,-1,-2,0,-1,-1,2,-1,1,1,0,0,-1,0,1,-1,-1,0,3,0,-1,0,1,1,-3,3,3,0,1,-1,0,0,0,-3,0,1,0,0,0,1};
			215: counter1_out = '{0,0,-1,0,0,2,-1,1,-1,-1,2,1,1,0,-1,-1,1,0,1,-2,0,1,0,0,1,2,0,2,1,0,0,-2,-2,0,0,-1,0,-2,0,0,0,0,-1,0,0,0,1,-1,-1,0,0,-1,0,1,0,0,2,-1,0,-1,2,0,-1,0,0,-1,2,0,1,0,1,0,-1,0,0,1,1,2,0,2,0,0,1,0,1,0,1,0,-2,0,0,1,0,0,-1,-2,1,-2,0,-1};
			216: counter1_out = '{1,-2,-1,1,1,2,2,1,2,1,1,0,0,1,1,0,0,-1,0,-1,1,1,1,1,1,0,2,0,0,0,0,0,-2,2,-1,1,1,1,-1,0,1,-1,0,1,-1,0,1,-1,0,1,0,1,1,0,-2,1,0,0,0,2,-1,-1,-2,1,1,-1,2,-2,0,1,0,-1,1,0,-1,0,1,2,-1,0,0,0,1,0,0,1,2,-1,-1,2,1,-1,1,-1,-1,1,-1,1,1,-1};
			217: counter1_out = '{0,1,0,1,0,2,0,1,-1,0,1,0,1,-2,0,0,1,1,-1,-1,0,-1,0,-1,-1,2,-2,1,0,2,1,-1,-1,0,2,0,0,-1,0,0,1,1,1,0,1,0,2,-1,0,1,0,0,0,-1,0,-1,-1,-1,0,1,0,-2,1,0,1,-1,1,-2,0,-1,0,-3,0,-1,0,0,0,1,-1,0,-2,-1,1,2,-1,-1,-1,0,0,1,0,0,0,-2,-2,0,-1,1,-1,1};
			218: counter1_out = '{1,-1,-2,0,1,0,2,0,0,0,2,1,0,0,-1,1,-2,0,0,-2,1,-1,0,1,-1,1,1,2,2,0,1,2,1,1,-1,-1,-2,2,1,-2,1,-1,-1,1,2,0,0,1,-1,-1,1,2,0,1,0,0,0,-1,0,0,-2,-1,0,0,1,1,1,0,1,1,-1,1,0,0,0,1,0,-1,0,1,2,-1,0,-1,-4,0,1,-1,0,2,0,-2,2,1,1,-1,-2,-1,0,-1};
			219: counter1_out = '{0,1,0,0,0,0,1,-1,-2,1,1,0,0,0,0,-1,2,1,-1,0,0,0,1,0,1,1,0,0,0,1,1,0,-1,0,0,1,-1,0,2,1,-1,0,0,-2,-1,-1,0,0,-1,1,1,2,3,2,2,0,-1,-1,0,0,0,0,-1,-2,-2,-2,0,1,-1,0,0,-1,0,0,-1,0,1,0,-1,1,0,1,0,-1,1,0,1,-2,1,2,1,1,1,0,0,-1,-1,0,1,-2};
			220: counter1_out = '{2,0,-1,-1,1,-2,-1,-2,1,0,0,1,0,1,-2,0,-1,1,-1,-1,1,0,-3,0,-1,1,-2,0,2,0,0,0,-1,-1,0,-1,1,-1,-1,0,2,0,0,0,1,-1,-1,0,-1,1,-1,0,0,0,0,-1,0,1,-1,-1,0,-1,0,-1,2,-2,1,-1,1,1,1,0,1,1,0,2,0,-1,-2,-1,-1,0,-1,0,2,2,0,-1,-1,0,1,-1,1,1,2,0,-1,0,1,-1};
			221: counter1_out = '{0,0,-1,0,0,2,-1,0,1,-1,0,0,0,2,-1,-1,-2,0,1,0,1,-1,0,0,0,1,0,0,1,-1,1,-2,-1,1,-1,-1,0,2,1,0,0,-1,-1,0,0,-1,2,-1,1,0,-1,1,0,0,0,2,0,0,-1,0,-1,1,2,-1,0,0,1,-1,1,0,0,0,0,1,-1,0,0,-1,0,0,-1,1,0,0,0,-1,0,1,-1,0,1,0,-1,0,-1,1,-1,0,-1,0};
			222: counter1_out = '{1,1,-1,2,1,-1,0,0,-1,1,0,1,2,-2,-1,-1,-1,0,0,0,1,0,-1,0,2,2,1,-2,0,-1,0,1,-1,-1,2,0,1,-2,-1,1,-2,0,0,0,0,1,0,0,-1,1,-1,0,2,0,1,-2,0,0,-1,-2,-1,1,2,-2,-1,1,1,1,-1,-1,0,1,0,1,0,-1,0,0,1,0,1,-1,0,0,-1,-1,-1,-1,-1,1,0,0,-1,-1,-1,0,0,1,0,3};
			223: counter1_out = '{-1,1,0,0,1,0,-1,0,1,0,0,1,1,-1,0,-1,-1,0,0,-2,0,0,0,0,-2,2,0,1,1,0,0,1,-1,-2,-1,1,0,1,-1,0,1,1,-1,1,-1,1,0,1,0,0,-1,0,0,-2,1,1,0,0,-1,0,1,1,0,-1,0,0,2,1,-1,2,0,1,-2,0,-1,0,1,-1,0,1,1,0,0,1,-1,0,0,-3,-1,-1,0,1,1,0,2,-1,-1,-1,-1,-1};
			224: counter1_out = '{1,0,0,1,1,1,0,-1,0,0,2,0,0,-1,0,-1,1,-2,0,0,0,-1,-1,0,2,1,1,0,-1,0,-1,0,-1,-1,0,-2,0,1,0,0,0,0,-1,-1,1,2,1,0,0,0,0,0,-2,1,0,0,2,1,2,-1,1,-1,0,-1,-1,2,1,2,0,-1,0,-1,-2,-1,-1,1,1,-2,2,1,0,0,-1,1,-1,1,0,1,1,-1,-1,1,-2,0,3,0,0,1,-1,1};
			225: counter1_out = '{1,1,-2,2,-1,0,1,1,0,0,0,-1,-1,1,0,-1,0,2,-1,-1,0,-1,0,1,-1,1,-1,0,0,-1,2,1,-1,0,0,0,1,1,0,2,-3,1,0,-2,-1,1,-2,-1,-2,-1,1,1,0,1,3,-1,-1,0,-1,-1,1,3,0,0,1,-1,0,0,1,3,1,1,1,-1,0,1,0,1,0,0,0,0,0,0,1,-1,1,1,-1,-1,-1,1,-2,-1,1,0,-1,-1,1,0};
			226: counter1_out = '{-1,-1,1,-2,-2,1,1,-1,0,-2,1,0,1,-1,-1,-1,0,-2,-1,1,0,1,1,0,1,1,-1,0,0,1,0,3,0,-1,-2,-1,2,0,-1,2,-1,1,-1,-1,-1,1,0,1,1,0,-1,-1,0,1,1,0,-1,0,0,-2,1,0,-2,-1,2,1,-1,2,-1,0,0,-2,-2,0,0,0,-1,-1,0,1,-1,1,-1,0,1,1,-1,-1,0,-1,0,0,1,-1,1,0,1,0,-1,0};
			227: counter1_out = '{2,0,-2,1,0,2,1,1,-1,-1,1,0,-1,1,0,0,0,1,-2,-1,1,0,1,-1,-1,1,-1,0,1,-1,-1,-1,2,1,0,0,-2,0,1,1,0,0,-1,-1,1,0,-1,-1,-1,0,2,0,0,0,0,0,1,1,0,1,1,0,0,0,-1,-1,0,1,1,1,0,0,0,-1,2,1,-1,1,2,2,0,1,0,-2,-2,0,1,0,0,0,0,-2,0,2,-1,2,0,0,-1,1};
			228: counter1_out = '{1,1,0,1,0,-1,0,1,0,1,0,-1,1,1,-1,0,1,1,1,-1,0,0,0,0,-1,2,1,0,0,1,1,0,1,-1,2,-1,-1,1,-2,-1,0,0,0,-1,0,0,-1,0,3,1,2,-2,1,0,-2,0,0,0,0,0,0,0,1,0,-1,-1,0,1,0,-1,0,1,-1,0,0,0,1,0,1,0,1,0,-2,1,0,0,-2,1,0,0,1,0,1,-2,-1,0,1,0,0,-1};
			229: counter1_out = '{0,1,-1,0,0,1,1,1,1,1,0,-1,-1,-1,2,0,0,1,1,-1,1,1,0,0,-1,-4,0,0,1,-1,0,-3,-1,0,2,1,-1,1,-1,2,1,1,-1,-2,-1,0,1,-2,-1,2,0,2,1,1,-1,1,-1,0,1,-1,0,-1,0,0,0,-1,-1,1,2,-1,1,0,0,0,1,0,1,2,-1,-1,0,0,1,0,-1,1,2,-2,-2,0,1,0,-1,1,0,0,-1,-1,0,0};
			230: counter1_out = '{1,-2,0,-1,1,0,0,0,0,0,2,0,-2,-1,0,-2,1,0,-1,-1,0,0,0,1,-1,1,0,-1,-1,0,2,1,0,0,0,1,-1,0,0,-1,0,0,-1,1,1,0,0,1,-1,-1,1,-2,1,1,-1,-1,0,0,0,1,-1,0,1,0,-1,1,0,0,1,0,0,1,-1,0,1,-1,0,1,0,-2,-1,-1,1,0,0,0,1,-1,-1,0,-1,0,-1,-2,1,2,0,1,-2,2};
			231: counter1_out = '{0,-1,0,0,0,0,0,0,2,0,-1,0,0,0,-2,1,-1,-1,-1,0,2,0,1,0,-1,1,-1,1,0,0,0,0,0,-1,-1,-1,-1,1,1,-1,-2,1,-1,-1,0,-2,-1,1,1,-1,0,-1,-1,0,1,0,1,0,1,-1,-2,0,-1,-1,0,1,0,1,0,-2,1,-1,1,1,1,1,0,0,0,0,0,-2,1,0,1,-1,0,0,-1,-2,0,0,-1,0,1,1,0,0,-1,0};
			232: counter1_out = '{0,-1,0,0,-1,1,1,1,1,2,-1,-1,1,-1,-1,-1,0,0,1,0,-1,1,-1,2,-1,0,1,0,0,0,-2,-1,2,-1,2,1,1,1,4,1,0,1,-2,-1,-1,0,-1,-1,1,-1,1,0,-1,1,-1,0,1,0,1,2,-2,-2,0,-1,0,1,1,0,1,0,-2,0,1,0,-1,0,-1,-2,1,0,1,0,0,-1,1,1,0,-1,1,-1,1,-1,1,-3,2,0,1,0,1,-1};
			233: counter1_out = '{-2,0,0,-1,0,0,0,0,0,-1,0,0,-2,1,-1,0,0,2,1,2,2,0,0,0,2,-1,1,-1,1,-1,0,-2,1,1,0,1,1,-1,1,-2,0,0,-1,0,-1,2,1,0,-1,-1,0,0,1,1,-1,0,0,0,-2,0,2,-1,0,1,2,2,1,-1,2,1,2,0,2,2,-1,0,0,0,0,0,0,1,1,1,-1,0,1,1,1,0,1,0,0,0,-1,1,-1,3,-1,2};
			234: counter1_out = '{0,-1,0,0,1,-1,-1,-2,0,2,-1,1,0,1,0,0,2,1,0,1,0,0,0,1,0,1,0,0,0,2,-1,0,0,-1,2,-2,-1,-2,-1,-1,0,0,1,0,1,1,0,0,1,-1,0,0,0,-1,2,2,1,2,1,1,-1,-1,0,-2,0,0,0,-1,0,0,1,-1,-1,0,1,-1,1,2,0,2,0,0,2,-2,-2,0,2,-3,-1,0,0,0,2,-1,1,-1,3,2,0,2};
			235: counter1_out = '{0,-1,-2,-1,-1,0,-1,-1,1,0,-1,2,-1,1,0,0,0,0,1,0,2,0,1,0,0,-1,0,-2,0,-1,-1,0,0,1,-1,-1,1,0,-3,1,-1,-3,-1,1,-1,0,0,-1,-1,-1,-1,0,0,1,0,-1,-1,-2,0,0,-1,-2,1,-1,-2,1,0,-2,0,-2,-1,-2,-1,0,-1,1,2,-2,1,-1,0,-2,1,0,1,0,3,-1,0,0,0,0,-1,0,-1,0,0,1,-1,-2};
			236: counter1_out = '{-1,0,-1,0,1,2,0,0,-1,0,0,2,0,-1,0,0,1,-1,2,0,-1,0,0,0,-1,0,0,-3,0,0,-1,2,-1,1,0,-2,0,0,0,1,-1,-2,0,0,-2,2,1,-1,0,1,-1,0,-2,0,-1,0,1,0,0,-1,1,-1,2,1,0,-2,0,0,2,0,2,-1,1,1,0,1,-2,0,-1,0,1,-1,1,-1,0,0,1,-1,-1,-1,0,0,-1,-1,1,0,-1,4,1,0};
			237: counter1_out = '{0,0,-2,1,1,1,2,0,-1,-1,1,-1,0,1,-1,-1,1,-2,1,0,-2,0,1,-1,0,1,0,1,0,0,-1,2,-2,0,1,2,0,1,0,0,-2,-1,0,0,0,0,-2,0,0,-1,-1,0,-1,-1,-1,-2,1,1,0,1,0,-1,2,-1,0,1,-1,0,-2,0,1,-1,0,-1,-3,0,0,1,0,0,-1,-2,1,1,0,-1,2,-1,0,2,1,1,1,0,0,0,1,2,0,0};
			238: counter1_out = '{2,1,1,1,0,4,2,1,0,0,1,1,-1,1,0,-1,1,-2,0,-2,0,-1,-1,-1,-2,-1,-1,-1,-1,-1,0,0,-1,-1,0,0,-1,0,-1,0,1,0,0,0,0,0,-2,-2,0,0,1,1,-1,-1,-1,-3,-4,1,2,-1,1,-1,2,-1,-1,0,0,-1,0,0,-1,0,1,0,0,-2,0,-1,-1,-1,0,1,0,-2,0,2,1,1,-1,0,-2,1,0,-1,0,-3,-1,2,0,-2};
			239: counter1_out = '{0,0,-1,0,1,3,-1,0,0,1,2,-1,-2,0,1,-1,-1,-1,0,1,1,1,1,-1,1,0,-1,-2,1,-1,1,1,-1,0,-2,-1,-1,0,1,1,0,-1,0,0,1,0,1,0,0,-1,3,0,0,-1,-1,-1,-2,-1,0,0,1,-2,-2,0,2,0,0,0,0,0,2,0,2,-1,1,-1,1,-1,0,0,-1,2,2,-1,0,0,4,0,0,-2,1,0,-2,0,0,-1,1,2,0,1};
			240: counter1_out = '{2,2,-1,1,0,4,-1,2,0,0,3,1,1,0,0,1,0,0,0,1,0,1,2,-1,-1,1,-1,0,0,0,0,0,-2,0,-1,-1,-2,-1,0,0,1,1,-1,0,1,1,0,-1,1,-1,3,0,1,-2,2,0,1,-1,0,0,0,-1,-1,-1,-2,0,-1,-1,-2,2,-1,-2,0,0,1,-1,1,0,0,0,-2,1,-1,-2,-2,0,1,0,0,0,1,-1,0,-1,1,-1,1,1,1,4};
			241: counter1_out = '{0,-2,-1,-1,1,2,-3,-2,0,1,1,0,0,0,2,0,-1,1,0,-1,0,0,0,-1,1,1,0,1,-1,0,0,-1,-1,-1,0,0,2,1,0,0,1,0,0,0,0,1,1,0,1,0,-1,1,1,0,1,0,1,-1,1,0,0,-1,-1,1,1,-1,0,-1,0,1,-1,-2,-1,-1,2,1,-1,1,1,1,-1,-1,1,0,1,-1,1,2,-2,1,-2,0,-1,-1,-1,-1,0,0,-1,3};
			242: counter1_out = '{0,0,-1,0,0,0,-1,0,0,0,2,1,2,1,0,1,0,-1,-1,0,1,0,1,2,2,1,2,1,0,0,0,-3,0,1,-2,-1,1,-1,-1,-1,0,0,-1,-1,0,1,0,-3,1,-1,2,2,2,-2,0,0,2,1,0,0,-3,0,-1,1,0,1,1,-1,-1,-2,0,-1,-4,-1,-1,0,-1,0,1,1,-1,1,0,-3,0,0,-1,0,0,-1,1,0,1,-1,1,1,1,-1,0,1};
			243: counter1_out = '{2,1,-1,1,1,2,0,-1,0,1,3,-1,0,0,-1,1,0,1,-1,0,3,0,0,-1,0,0,0,-1,-1,0,1,0,-2,0,2,-2,0,2,-2,-2,-2,-1,-1,1,-1,0,1,0,0,-1,1,0,0,-1,2,0,0,0,0,0,0,0,0,0,-1,0,3,0,-1,0,0,0,-1,-2,-2,1,1,-1,-1,0,0,-2,1,0,-2,0,0,-1,-2,1,0,0,1,-2,-1,0,0,0,0,0};
			244: counter1_out = '{-3,1,-2,1,-1,0,1,0,1,0,3,1,0,1,-2,1,0,0,-1,1,-1,0,1,-1,-1,0,0,0,-1,0,-1,0,-1,-1,0,2,0,-1,1,1,0,0,0,0,1,1,-2,-1,-1,1,1,2,0,0,-1,-1,1,0,1,0,1,-2,-1,-1,0,1,1,0,0,0,1,2,-2,0,-1,2,-1,0,2,1,0,0,1,-1,1,2,0,-1,2,0,0,-1,0,0,0,-1,-1,0,0,0};
			245: counter1_out = '{-2,1,-1,-1,2,2,1,0,1,-1,1,1,-1,0,0,-2,1,-1,-2,0,1,-1,-1,1,0,0,1,2,-1,-1,0,0,0,0,0,1,0,2,0,0,0,0,-1,0,0,0,-1,-1,-3,1,0,-2,0,-2,-1,1,0,-2,1,0,1,0,0,1,0,0,1,0,-1,0,0,1,-1,1,0,-2,2,1,-1,0,1,1,1,0,-1,-1,1,0,-2,0,0,0,1,-2,0,-2,1,-1,1,-1};
			246: counter1_out = '{0,0,-1,1,0,0,0,1,-2,1,3,1,-1,-1,1,-1,0,1,-1,0,-1,-2,0,0,-1,0,1,-1,0,0,2,0,-2,0,0,-1,-1,-1,1,0,-1,1,0,0,0,1,1,-4,-1,-1,0,0,1,-1,0,1,0,0,0,0,0,0,-3,-1,-1,-2,0,0,-2,-1,0,1,1,1,-1,1,2,-2,1,0,-1,1,2,1,1,1,0,0,-2,2,1,1,2,-1,0,0,-1,-2,-2,0};
			247: counter1_out = '{1,2,0,0,1,1,1,1,0,0,1,-1,0,-1,0,-2,2,1,-1,-1,0,1,0,0,2,1,1,-1,-2,1,1,1,1,-1,0,0,-2,1,2,1,-1,-1,-1,-1,0,1,-1,1,-3,0,-1,1,-1,-1,2,-1,1,-1,1,0,-2,0,-1,-1,-1,-1,0,-1,0,0,0,1,1,-1,-1,2,2,1,-1,0,-2,1,3,1,1,0,0,1,-2,2,0,0,0,0,1,0,-2,1,1,-1};
			248: counter1_out = '{1,-1,0,-1,0,-2,0,0,0,1,1,0,1,0,0,-1,0,0,0,-1,-1,1,-1,0,-1,1,1,2,0,-1,-1,1,-1,0,0,0,-2,2,1,1,-1,1,0,-1,1,-1,-1,0,-1,1,-1,1,0,1,1,0,3,1,-1,-1,0,0,0,-1,0,0,1,0,-1,0,-1,-1,0,0,-1,1,-1,-1,1,0,1,1,1,1,0,-1,0,0,0,1,0,-1,0,1,0,1,-2,2,-1,2};
			249: counter1_out = '{1,0,2,1,-1,0,2,1,2,1,-1,-1,0,1,1,-1,0,0,-2,0,0,0,-2,-1,1,1,0,1,1,-1,-1,0,0,0,1,-2,1,1,0,-1,0,1,1,-1,1,-2,0,0,1,0,2,-2,-1,0,2,0,-1,1,0,-1,0,1,-1,0,0,0,0,0,1,1,1,-2,-4,1,-2,0,1,1,-1,-2,0,0,1,-1,0,2,0,-1,-1,-1,-1,0,-1,0,0,-1,-1,1,-1,-1};
			250: counter1_out = '{0,-1,-1,0,0,-1,2,0,0,-1,1,0,0,0,-1,-1,0,2,0,-1,-2,-2,0,-1,-2,-2,-1,-1,0,-1,1,-1,2,2,0,0,0,0,0,0,1,1,0,0,0,-1,-1,1,0,0,2,-2,1,1,0,0,-1,1,1,0,1,-1,0,1,-1,0,0,0,1,0,1,1,1,0,-1,1,1,0,0,0,-2,-2,0,1,1,-2,2,0,-1,0,-1,-1,0,1,-1,0,0,0,1,1};
			251: counter1_out = '{0,0,1,1,1,0,1,0,0,0,1,1,1,0,0,1,0,0,1,0,-4,-1,-1,0,0,-1,-1,2,0,1,0,2,0,-1,0,0,0,0,0,0,-2,0,0,1,0,-1,-1,2,0,0,0,-1,-3,2,0,0,0,0,1,0,-1,1,0,0,1,1,0,0,-1,0,0,0,1,1,1,1,-1,2,0,0,1,0,1,-2,0,-1,0,0,-1,-1,0,-1,0,2,1,0,0,-3,0,1};
			252: counter1_out = '{2,0,-1,0,1,2,-2,0,0,-1,2,0,-1,-1,0,-1,1,0,0,0,-1,-1,-2,1,1,1,0,0,2,0,-1,0,0,0,1,-1,-1,1,-1,-1,1,0,0,-1,1,0,-1,-1,1,0,-1,1,-1,1,1,0,-1,0,-2,0,3,1,0,0,0,-1,1,-1,0,1,-1,0,1,1,2,-1,-1,1,0,0,-2,-2,0,-1,-1,-1,-2,2,1,0,2,0,0,1,0,0,0,-1,1,-1};
			253: counter1_out = '{1,1,0,-2,-1,-1,2,0,-2,0,-1,0,-2,1,-1,-1,1,2,-1,-1,-1,1,0,0,1,0,2,-1,1,0,0,-1,2,-1,0,0,0,-1,1,-1,-1,-2,0,0,-2,1,0,1,0,-2,0,1,1,-1,0,1,0,0,-1,-2,-1,0,0,-1,0,0,-1,0,0,0,1,2,1,-1,1,0,0,0,-1,-1,-3,0,2,0,-1,1,-1,-2,1,1,0,0,0,-1,0,0,-2,1,0,0};
			254: counter1_out = '{0,-1,1,-1,1,-1,0,-1,-1,0,-1,0,0,-1,0,2,1,0,0,-1,-1,-1,1,0,1,1,-1,2,0,-1,2,0,-1,0,1,1,-1,0,-1,1,0,1,-1,0,-1,1,1,1,1,2,0,-1,0,0,1,1,0,1,0,0,-1,0,0,1,0,2,0,0,-1,-1,0,1,-1,1,1,0,0,1,-1,0,1,0,1,-1,-1,-3,0,1,1,-1,-1,-1,0,0,-1,1,2,1,-3,1};
			255: counter1_out = '{-2,1,0,0,0,1,0,0,1,0,-1,-1,-1,1,0,0,0,0,0,-1,-1,1,-1,0,0,0,1,0,0,-1,1,1,-1,0,0,-2,-1,0,1,0,-3,-1,1,2,1,1,-1,1,-1,-1,1,0,2,0,0,0,-2,2,1,0,0,-1,0,1,1,1,-1,1,1,2,0,-1,1,-1,1,1,1,-1,0,1,-1,-2,1,0,-1,1,-1,0,2,-1,0,1,0,-2,0,-1,2,0,0,-1};
			256: counter1_out = '{0,1,-1,0,-1,0,-1,2,-1,1,1,-1,1,0,1,0,1,-1,0,0,-1,0,0,1,0,0,-1,0,1,2,2,0,0,1,1,1,-2,0,2,0,1,0,-2,0,-1,0,1,1,-1,2,1,0,0,1,-1,-1,0,-1,-1,-1,-1,0,1,2,0,0,1,0,0,0,1,0,1,1,1,0,-1,0,0,0,0,0,2,-1,0,1,0,0,-1,0,0,2,1,1,1,0,-1,0,-1,2};
			257: counter1_out = '{0,0,-1,0,0,-1,0,-1,-1,-1,2,0,1,0,-1,-1,0,0,1,1,0,0,0,1,1,-1,1,0,1,-1,-1,-1,1,3,1,1,2,-2,0,0,0,1,0,-2,1,-2,1,-1,0,0,0,1,0,0,0,2,-1,0,-1,1,1,1,-1,1,-2,0,-1,0,0,0,1,-2,2,0,1,3,2,-1,1,0,0,-1,-1,3,0,0,-1,1,0,1,0,-2,2,-1,1,-2,-1,-2,0,0};
			258: counter1_out = '{1,0,0,-2,-1,0,-1,0,0,2,0,2,0,1,-1,0,3,1,0,2,1,0,0,1,1,0,-3,-2,0,-1,0,-1,0,0,0,-1,0,0,0,0,0,-2,-1,-1,0,1,0,1,2,0,0,0,-1,1,1,-2,-1,0,-2,0,1,-1,0,-2,2,1,1,0,2,0,2,0,-1,-2,-2,-1,2,1,2,0,1,0,2,2,0,2,1,2,1,1,-1,-1,0,-2,1,-1,1,-1,0,1};
			259: counter1_out = '{0,-1,-1,0,1,-1,-1,0,1,0,-1,0,1,1,0,1,1,-1,-1,1,-1,0,-1,0,0,-1,0,0,0,1,2,-2,1,0,0,-1,-2,-1,1,-1,1,0,0,0,-2,0,1,-1,0,2,-1,1,-3,0,0,-2,1,1,-1,1,2,-1,-1,0,2,0,-2,-1,0,1,2,0,-2,-1,-1,0,-1,1,0,0,0,-1,0,0,-1,1,1,1,-2,-1,-1,0,1,-2,0,0,0,0,0,1};
			260: counter1_out = '{-1,-1,0,-2,-1,-1,0,0,-1,1,-1,-1,1,-1,1,-1,-1,1,-1,0,1,0,-1,-1,-1,-1,0,-1,0,-1,0,0,1,-2,1,0,0,0,2,1,0,1,1,-1,-1,2,1,-1,-1,1,0,-1,0,-1,0,-2,-2,1,-1,-1,-1,1,2,0,1,-2,1,0,-1,-1,0,1,0,-1,-2,1,2,0,-1,-1,-1,1,-1,-1,0,2,-1,1,-1,0,0,0,-1,-2,1,0,-1,1,-1,0};
			261: counter1_out = '{0,-1,1,-2,0,1,-1,0,-1,1,0,-1,-1,-1,-1,-2,0,1,1,1,-1,1,0,1,2,-1,-1,-2,-1,-1,0,1,0,-2,1,1,-1,-1,1,-1,-1,0,-1,-1,1,0,0,-1,-2,0,-2,1,-1,-1,-2,0,-1,-1,0,0,0,-2,0,2,1,-1,-1,-1,1,0,1,0,1,2,0,-2,1,1,1,-1,-1,-2,0,0,0,-1,1,-1,0,-1,3,2,1,0,0,1,-2,1,-1,1};
			262: counter1_out = '{-2,-3,-2,2,0,1,2,0,-1,0,-1,0,1,-1,1,-1,0,1,0,0,0,1,0,-2,0,0,0,0,0,-1,-1,0,-2,1,-1,-1,2,0,0,2,0,-1,-2,1,1,0,0,0,-1,1,0,0,1,0,-1,2,0,0,-2,0,2,-1,-1,-2,-1,-1,0,0,1,-1,3,1,-2,0,-1,1,0,0,0,-1,-1,0,-1,-1,-1,1,1,0,-2,0,-1,0,0,-2,0,0,-1,2,-1,-1};
			263: counter1_out = '{0,-1,-1,1,-1,0,-1,-1,1,-1,0,0,-1,2,0,-1,0,1,-1,-1,0,0,-1,-2,-1,1,-1,0,0,-1,1,1,0,1,0,1,0,0,0,1,-2,0,-1,0,-3,2,-1,-2,-2,1,0,-2,1,0,-1,0,0,1,1,1,1,-1,1,0,0,0,0,-2,-2,1,2,2,-2,-1,-2,1,1,0,0,-1,-1,-2,1,-3,-2,-1,0,-2,-1,-1,-1,-1,1,-2,1,2,-1,0,1,0};
			264: counter1_out = '{-2,-2,1,0,1,0,1,1,0,0,2,0,0,0,-1,-1,-1,1,-1,0,0,1,0,-2,2,-1,0,-1,1,0,-1,-1,-3,-1,1,0,1,0,-1,2,-1,0,-2,1,-1,1,-2,-1,-1,0,-2,0,-2,0,0,1,0,1,2,-1,2,-1,0,-2,1,-1,1,-2,0,0,2,2,-1,1,-2,0,-1,-1,0,0,0,-2,2,-1,1,0,0,-2,-1,-1,0,2,3,0,0,0,0,0,-1,0};
			265: counter1_out = '{1,2,-2,-1,0,0,0,1,-2,0,1,-1,-1,-1,3,-2,-1,-3,0,2,0,-2,-1,0,0,1,0,-1,1,-1,1,1,0,1,1,-2,1,1,-1,-2,0,-1,-1,0,-1,2,-1,-1,0,0,1,1,-1,0,1,-1,-2,1,0,0,1,-1,1,1,-2,1,-1,0,0,1,4,2,2,1,-2,0,2,-1,-1,-2,0,-1,1,1,-3,-1,0,1,0,-1,1,1,0,0,1,-1,2,-3,-1,-1};
			266: counter1_out = '{0,1,0,-1,0,-1,1,1,0,2,2,0,1,-1,1,0,-1,-1,1,1,-1,0,-3,0,0,-2,0,-2,-1,-1,0,0,-2,0,0,2,-1,0,0,-1,1,-2,0,1,-1,2,-1,0,0,-1,1,-2,0,2,0,-2,0,-1,0,1,0,-2,1,0,0,-1,-3,0,-2,1,3,-1,1,1,-1,1,0,1,0,-2,-1,-1,2,-1,-2,2,2,3,1,0,-3,0,1,-1,0,-1,1,-2,-1,1};
			267: counter1_out = '{0,0,0,0,0,0,-1,1,-1,1,1,-2,1,-3,1,0,-2,0,-1,2,0,0,-2,-3,1,-1,-1,1,-1,-1,-1,-1,-1,1,-1,0,0,1,2,0,1,0,1,0,-1,1,-1,-1,0,1,1,0,1,0,1,-2,-2,-3,1,-1,-1,-3,0,-1,-1,1,-2,-2,-2,-1,-1,0,1,-1,1,-1,-1,1,1,0,1,1,1,1,-1,1,1,2,0,-1,-2,-1,1,-1,0,1,2,0,1,3};
			268: counter1_out = '{1,-1,0,0,1,2,0,1,-2,-1,4,0,1,0,1,0,0,2,-2,1,1,0,1,0,1,-2,0,-2,0,-1,1,-1,-1,1,0,-1,1,-1,0,0,1,-1,1,0,1,0,2,-1,0,-1,1,1,1,1,0,1,0,0,1,-1,-3,-1,-2,0,0,1,-3,0,-2,0,0,-1,-1,-1,-1,-1,1,-1,2,-1,0,-1,2,0,-1,-1,-1,1,0,-1,1,0,0,-1,0,0,1,-3,-1,5};
			269: counter1_out = '{-2,1,0,1,0,1,-2,0,0,1,3,-1,0,-1,0,-1,-1,1,1,2,3,2,1,-1,1,0,-2,-2,1,1,0,1,0,2,1,1,2,2,1,0,0,1,0,-2,-1,0,0,1,1,0,1,1,0,-1,-1,0,0,-2,0,-1,1,-2,-2,2,-1,1,3,0,0,-2,1,0,0,1,0,0,0,1,-1,0,0,2,1,1,-1,0,0,-1,-1,-1,0,-1,2,-1,1,-1,-1,1,0,0};
			270: counter1_out = '{-1,0,-1,0,1,2,0,1,-1,0,0,-1,3,0,0,2,2,1,-2,0,0,-1,-1,0,1,-2,0,-3,0,2,1,1,-1,3,0,0,1,1,3,0,0,-1,0,-1,1,-1,1,0,0,0,1,1,2,-1,1,0,-2,-5,1,0,1,-2,0,0,0,-1,4,1,-2,-2,0,1,1,0,1,1,1,-1,0,2,1,1,1,0,-2,0,0,-1,-2,-1,1,-1,1,-1,1,0,1,0,0,-2};
			271: counter1_out = '{0,0,0,0,1,2,-1,1,-1,0,1,0,-3,-1,-1,0,-1,-2,-1,1,1,0,0,0,0,-3,2,-2,0,0,-1,0,2,-1,-1,-1,1,0,1,0,-2,1,0,-2,-1,1,1,0,0,0,0,0,1,-1,2,1,2,-1,0,-1,-1,1,-1,-1,1,1,2,-1,0,-1,-1,-2,-1,0,0,-1,0,0,0,0,-1,0,1,1,-1,0,0,-1,0,-1,-1,-2,0,0,2,0,2,1,2,-1};
			272: counter1_out = '{1,1,-1,0,0,-1,3,1,1,0,2,0,0,-1,2,2,1,0,-1,-1,0,0,-1,-1,0,-1,1,0,0,1,0,0,-1,1,0,1,2,1,1,-1,-1,-1,-1,-2,1,-1,-1,0,-1,-2,1,0,0,2,-1,1,-1,-2,1,1,0,0,-1,3,-1,0,2,2,-1,0,0,0,0,0,-1,1,1,0,1,1,1,-1,0,-1,-1,0,2,-1,2,0,0,1,0,0,0,-1,0,-1,0,-1};
			273: counter1_out = '{-2,0,0,0,-1,0,2,-1,0,0,0,-1,-1,-1,0,0,2,-1,1,0,0,0,0,1,1,-1,-1,0,0,1,0,0,-1,-1,1,0,0,2,1,-1,0,-1,0,-2,-1,-1,-1,1,-3,0,0,-1,-2,1,-1,-1,1,-4,0,-1,-1,1,0,1,-1,0,2,2,-1,0,1,1,1,1,-1,0,0,0,1,1,-1,0,-1,1,-1,0,-2,-1,-1,-3,1,0,1,1,2,0,0,-2,0,0};
			274: counter1_out = '{1,1,1,1,-1,1,0,-1,0,2,2,-2,0,-1,0,-1,0,-1,0,1,0,1,0,-1,1,-2,0,-1,-1,1,2,0,0,0,1,-2,0,0,0,2,-2,0,0,-2,-2,1,-1,1,-1,0,1,1,1,0,2,1,0,-3,2,1,0,1,-2,-3,1,0,1,2,-1,-1,0,1,0,-1,1,0,2,1,2,-1,-3,0,0,1,2,1,-1,0,-1,-1,1,0,0,1,2,1,1,0,2,-1};
			275: counter1_out = '{-2,0,0,0,0,-2,2,0,-2,1,1,-1,1,-1,-1,-2,-1,0,0,0,-3,-1,0,0,-1,0,0,-1,-2,0,1,-1,0,-1,-1,0,0,0,1,0,1,1,-1,-3,0,-2,1,-1,-1,-1,1,-1,0,0,1,-1,2,-1,1,1,1,-1,-1,1,-1,-1,0,2,-2,-1,2,0,0,-1,-1,-1,0,0,0,2,-1,0,0,1,0,-2,-2,-3,-2,0,1,1,1,-1,-1,-1,1,0,1,-1};
			276: counter1_out = '{-2,1,-1,1,-1,0,2,0,2,1,0,1,1,0,0,1,1,-1,-1,0,0,-1,-1,-2,1,0,0,0,1,0,-1,2,0,1,1,-2,-2,2,0,-1,1,1,1,-2,-1,-1,-2,1,0,-2,1,1,1,0,0,-1,0,-1,0,-1,-1,-1,-2,0,0,0,0,-1,1,0,-1,-1,0,-1,0,1,0,0,1,1,3,-1,-1,-1,1,-2,1,-1,0,-1,0,-2,1,-1,0,1,0,2,-1,0};
			277: counter1_out = '{-1,1,-1,0,-2,0,-1,0,-1,3,1,0,1,0,0,-1,1,0,1,0,-1,-1,-1,0,1,1,0,0,0,0,2,1,1,-2,-1,0,-2,-1,1,0,1,1,1,1,0,0,0,0,-1,-1,-1,1,-1,0,1,1,0,0,1,0,0,0,1,0,0,1,0,0,-1,-1,0,1,0,-1,-1,0,2,1,0,1,1,-1,1,1,-1,1,-1,-1,0,1,0,-1,1,0,0,-1,1,2,1,1};
			278: counter1_out = '{0,1,-2,-3,0,1,0,1,-2,1,0,1,0,1,-1,0,-1,1,-1,0,0,-1,0,2,-1,-1,0,2,0,0,0,1,0,0,0,1,1,-1,1,1,0,1,-1,0,0,1,0,1,0,-1,1,-1,2,-1,-2,0,0,1,-1,0,0,1,0,-1,0,1,0,1,0,-1,0,-2,-2,0,0,-1,-1,0,1,0,1,1,1,2,0,1,-2,-1,1,0,1,-2,0,0,-1,0,0,0,0,-1};
			279: counter1_out = '{0,1,0,0,1,0,2,2,-2,0,0,-2,0,1,-2,1,-1,0,0,0,1,0,0,0,-2,2,1,0,-1,-3,0,1,-1,-2,-1,2,-2,2,-1,-1,-2,-1,0,2,0,-2,0,0,2,-1,0,1,0,1,-1,1,1,-1,-1,0,1,0,-1,0,-1,1,0,0,1,0,0,-2,1,1,0,-1,-1,0,0,0,0,-1,1,-1,0,0,1,1,0,-1,1,0,0,0,0,-1,0,1,0,0};
			280: counter1_out = '{2,-1,-1,0,-1,1,1,0,2,1,-1,-1,-1,1,1,2,-2,-2,0,-2,1,-1,0,0,-1,-1,0,1,-1,0,-1,-1,0,-1,0,1,2,0,-1,-1,-1,1,0,0,-2,0,1,1,1,1,0,1,2,0,0,1,2,-2,-1,-1,1,0,2,0,-1,-1,1,0,2,-2,2,-1,1,1,2,-1,1,-1,-1,0,-1,-1,0,2,0,0,0,0,1,-1,0,0,-2,-1,-1,-1,0,1,0,2};
			281: counter1_out = '{0,1,0,0,0,-1,0,0,-2,1,0,1,-1,0,1,0,-2,-3,-1,0,1,-1,0,-1,0,1,0,0,1,1,0,0,-1,0,0,0,-1,-2,-1,0,1,0,-1,-2,0,1,2,1,-1,0,0,2,1,0,1,0,2,-2,0,0,-1,0,-1,2,1,0,1,0,0,2,-1,-1,1,1,0,-1,-1,1,-1,-1,1,-2,0,0,0,2,0,1,-1,1,1,1,0,-1,2,-1,-1,0,0,-1};
			282: counter1_out = '{0,0,1,-1,-1,1,-2,2,-1,0,-2,-1,-1,0,-3,0,1,0,-1,0,2,-1,-1,3,1,0,0,2,-2,-1,0,1,-3,1,0,0,0,1,0,0,0,0,-1,0,1,2,1,0,1,-2,1,0,0,2,0,1,2,1,3,-1,1,0,0,0,0,0,0,1,1,1,0,0,0,0,-1,0,-1,-1,-1,-1,1,-1,-2,0,1,1,-1,-1,1,2,0,-1,1,2,1,0,1,0,2,-1};
			283: counter1_out = '{1,-1,0,0,0,0,-1,0,1,0,1,0,-1,-1,-1,1,0,0,0,0,1,-1,-1,-1,1,0,-1,2,0,0,1,-2,0,1,2,1,1,0,0,1,1,1,0,1,-1,1,0,1,0,0,0,0,-1,1,-1,0,0,-2,2,1,1,-1,-1,0,0,0,0,0,2,1,0,1,-2,1,0,0,-1,0,1,-1,1,-1,2,1,1,-1,0,1,-2,0,-1,2,-1,0,0,0,0,-2,-1,-1};
			284: counter1_out = '{-2,0,-1,0,0,0,1,1,0,1,1,1,0,0,-1,1,-2,0,0,0,1,1,-1,2,0,0,-1,-2,-1,-1,0,1,0,-1,1,2,0,-1,0,-1,1,0,0,0,0,0,-1,0,2,0,-2,0,1,1,-2,-2,-1,0,-1,0,-1,-1,1,0,-1,-1,-1,0,0,-2,2,0,0,1,0,2,0,0,0,2,0,1,2,-1,0,1,-2,-1,-1,-1,0,0,-1,-2,-2,0,-3,-1,-1,1};
			285: counter1_out = '{-3,1,0,1,-1,0,0,-1,1,-1,2,-1,-1,-2,0,0,0,0,-1,0,0,-1,-1,2,0,1,0,1,-2,1,-2,1,1,-1,0,-2,0,0,-1,1,0,0,0,-2,1,1,-1,1,0,1,1,0,-1,-2,0,2,1,-1,1,1,0,0,-2,1,3,1,-1,0,-1,1,0,0,0,2,-2,-1,1,0,0,1,1,0,-2,-1,2,0,-1,-1,0,2,0,0,-1,0,1,0,-1,0,1,-1};
			286: counter1_out = '{1,-1,0,2,1,0,0,-1,3,-1,1,-1,-1,1,0,-2,2,0,1,0,0,0,0,-1,-1,-1,0,1,0,0,1,0,-2,1,-1,0,0,0,1,0,0,0,0,0,-1,2,-1,0,0,-1,0,0,1,-1,-2,-2,0,0,1,1,1,0,-1,-2,2,1,0,-2,1,0,2,0,0,0,0,2,1,-1,-1,1,0,-1,0,1,1,-1,1,-1,0,-2,-1,1,1,0,2,-1,-1,0,1,1};
			287: counter1_out = '{-1,0,0,-1,1,1,0,0,0,0,-1,0,0,0,-1,-1,0,1,1,-1,-2,0,-1,0,0,0,0,-1,-1,-1,1,-2,-1,-1,0,0,-1,1,2,1,1,0,1,-2,-1,0,0,-1,-1,0,0,-1,-1,-1,0,0,0,-2,-1,-2,0,0,-1,0,2,1,0,-2,0,0,-1,-1,2,0,-2,0,-1,1,-1,-1,0,0,1,-2,1,0,0,0,0,-1,-1,0,-1,-2,0,0,0,0,-1,1};
			288: counter1_out = '{0,0,1,-1,-1,-2,-1,1,-2,-1,0,1,0,2,-1,-2,2,1,1,1,1,0,0,1,1,0,-2,1,0,1,-1,0,-2,1,-1,1,0,1,2,-1,1,1,0,0,1,2,0,-1,-2,1,0,0,0,-1,-1,-1,0,1,0,0,0,1,-1,0,1,0,-1,1,0,0,0,0,0,0,-3,-1,3,0,1,-2,0,1,1,-1,1,0,0,-1,0,-2,-1,-2,0,-2,0,1,0,0,-1,0};
			289: counter1_out = '{0,1,2,-2,1,0,0,0,0,-1,0,0,0,0,1,-2,1,1,-1,0,-2,2,-2,0,0,1,1,-2,-1,0,-1,-2,-2,1,0,0,0,0,-2,0,1,0,0,-1,0,1,1,-1,-2,0,0,1,-1,-1,1,1,1,0,1,0,1,1,0,0,1,0,0,-2,1,-1,-1,1,-2,-1,-1,0,-2,0,2,-1,-2,-1,-2,0,1,-1,1,1,0,-1,1,-1,0,1,1,0,-1,-1,-1,0};
			290: counter1_out = '{-1,-1,-1,0,1,0,2,0,-1,-1,0,0,1,1,1,-2,1,1,-2,1,1,1,-4,0,-2,1,1,-1,0,0,-2,1,-1,-1,0,2,-1,0,1,-1,0,-1,0,-1,-1,0,0,0,-3,0,0,0,0,-2,1,0,0,0,1,-2,-1,0,-2,-1,-1,0,-1,1,0,0,1,1,-1,0,-3,0,1,-1,-2,0,1,-1,1,0,0,2,0,0,0,-1,1,0,0,0,0,-1,0,0,-1,1};
			291: counter1_out = '{1,0,-1,2,-1,-1,-1,1,0,-2,0,1,3,-3,0,-1,1,0,0,1,1,0,-4,0,0,-1,-1,-2,0,-1,0,1,-1,0,-2,-1,-1,0,-1,-2,-1,0,0,0,-1,1,-1,0,-2,0,-1,1,2,-1,1,2,0,0,0,0,0,-1,0,0,0,0,-2,-1,0,1,0,1,-2,0,-1,2,0,-1,2,-1,-1,0,-1,-2,0,0,-1,-1,0,2,2,-1,0,-1,1,2,-1,0,1,0};
			292: counter1_out = '{-3,-1,1,2,0,0,0,0,-1,-1,2,0,0,1,1,-1,0,0,0,0,-1,0,-3,0,-1,1,-1,1,0,0,0,0,0,0,0,-1,-1,0,0,1,0,0,0,0,0,1,-1,-3,0,0,-1,0,0,0,1,0,-2,0,0,-1,1,2,-1,0,1,0,-1,-1,0,-1,1,2,0,-1,0,3,1,1,1,-2,-1,-2,0,-1,1,0,1,0,0,0,1,2,0,0,1,-1,0,-3,2,-1};
			293: counter1_out = '{-2,0,-2,1,1,0,0,0,1,-1,0,-3,0,1,0,0,0,-3,1,0,-1,0,-3,0,-1,-1,0,-3,-2,0,2,-1,-1,2,2,0,-4,0,-2,0,1,-4,-2,-1,-1,2,-3,-1,2,-1,1,0,0,2,1,-4,-1,0,1,0,1,1,2,-1,-2,-1,-3,-1,-2,0,1,0,1,-1,-1,1,1,1,1,1,1,-4,4,0,1,0,1,2,-1,1,1,0,2,2,0,0,-1,-1,0,-1};
			294: counter1_out = '{-1,0,-3,-1,0,-1,0,0,1,-1,-1,-1,1,0,0,0,-2,-3,1,2,1,1,-3,0,-1,-1,0,0,0,-2,0,1,-2,1,-1,0,-3,1,0,2,1,-1,1,-1,0,3,-1,-1,2,-1,0,0,1,0,1,-1,0,-2,1,0,0,0,2,-1,0,0,-3,0,0,0,2,1,1,1,0,-1,0,0,0,-1,-2,-1,1,1,1,1,-1,0,-1,-1,1,-1,1,1,1,0,0,-3,0,2};
			295: counter1_out = '{1,0,-1,0,1,0,-1,0,1,1,2,-1,1,-1,1,1,-2,0,-1,1,1,0,-1,-1,1,-3,0,0,1,-1,1,0,1,-1,-1,0,0,0,-1,0,1,0,1,1,-1,1,-1,0,0,-1,3,0,1,-1,1,2,0,0,2,0,1,1,-3,-2,0,0,0,1,-2,0,-1,1,1,2,0,1,-1,0,1,0,1,1,1,-1,-1,-1,-1,3,-1,-1,0,0,1,0,-2,-1,1,0,-1,3};
			296: counter1_out = '{0,0,-1,1,0,-1,-1,0,-2,0,-1,-2,0,-2,1,2,2,0,-1,0,2,1,2,0,0,-3,-1,-3,-1,-2,1,0,1,1,-2,0,0,-1,0,1,-1,0,0,0,-1,1,2,1,0,0,2,-1,-1,1,1,0,1,-2,2,1,1,2,0,0,0,1,-1,0,-1,0,0,1,1,0,1,-1,1,0,-1,2,-1,2,2,1,-2,-1,-1,2,0,-1,0,-3,4,1,1,2,0,-2,0,1};
			297: counter1_out = '{-1,2,0,-1,0,-1,-2,1,1,1,1,-1,-1,-1,1,0,2,-1,-2,1,1,-1,0,0,1,-3,-2,-4,-1,-1,-1,-3,-1,-1,0,-3,3,-1,0,1,-1,0,1,-2,0,-1,1,0,1,-1,0,0,0,0,0,0,0,-2,1,0,1,1,0,0,0,1,-1,2,0,1,0,1,0,0,0,-1,-1,-1,0,1,2,-1,3,1,-2,2,0,-1,1,0,-2,-1,0,1,1,1,1,2,0,1};
			298: counter1_out = '{0,0,-1,2,0,0,2,0,-1,-1,0,-1,1,-3,0,0,-2,-1,0,2,0,2,1,1,-2,-2,-2,-1,-1,0,2,1,1,-1,0,2,1,0,1,2,0,0,0,-2,-3,1,1,2,0,0,1,0,0,1,1,0,0,-2,1,-1,1,1,-1,0,1,1,3,1,0,-1,0,1,-2,-1,0,-1,1,0,-1,-1,1,0,2,-1,-2,-1,0,-1,0,-1,1,2,-1,0,1,-2,1,-1,1,-2};
			299: counter1_out = '{-1,0,1,0,2,0,1,0,-1,0,-1,-2,0,-2,0,0,0,0,1,2,1,3,0,0,-1,-2,2,-1,1,1,1,-1,-1,0,0,0,0,-1,2,3,0,1,0,0,-1,0,1,2,-1,-1,1,1,0,1,0,-1,2,-4,1,1,1,-1,-1,1,0,1,1,3,-2,-1,1,1,-1,0,1,1,-1,0,-1,0,1,1,1,-2,-3,1,-1,-1,2,-1,-1,1,0,-1,0,2,1,1,-2,-2};
			300: counter1_out = '{-1,0,0,1,0,0,0,1,0,1,1,0,1,0,1,-2,0,0,2,1,0,0,1,0,0,-3,2,0,-1,2,0,1,1,-2,0,1,-1,1,1,0,-1,0,0,-2,-2,2,0,2,-2,-2,0,2,1,-3,-1,0,0,-3,-1,0,2,0,0,2,-2,0,1,1,0,-2,-2,0,0,1,1,0,1,0,-1,1,-2,-2,0,1,0,1,-1,-2,0,-2,1,1,0,0,2,0,1,0,0,-1};
			301: counter1_out = '{-2,2,0,1,-1,0,2,0,0,0,2,-3,1,-2,1,1,0,-1,-1,1,0,1,1,-1,0,-4,0,0,2,0,-1,2,-1,1,1,-1,-2,0,1,-1,2,0,-1,-1,-2,-1,-1,1,0,-2,-1,1,1,-1,-1,1,-1,-3,-1,1,-1,-2,-1,-1,-2,0,0,1,-2,-1,2,0,1,0,0,1,-1,1,1,0,0,1,1,-1,-2,0,-1,-1,-1,-1,1,-1,-2,-1,1,-2,1,2,0,0};
			302: counter1_out = '{0,2,1,2,3,1,1,2,0,-1,1,1,-1,-1,1,-2,1,1,0,0,-1,0,1,-1,-1,-1,1,-2,1,0,0,0,-1,-1,1,1,0,2,2,0,0,0,0,-1,0,-1,0,2,0,-1,-1,1,0,-2,0,-1,0,-1,0,-1,1,0,-1,-1,0,1,2,2,-1,2,0,0,1,2,0,-1,-1,1,0,0,-1,1,-1,0,1,0,-2,-1,0,-1,-1,3,1,1,2,2,3,0,0,-1};
			303: counter1_out = '{2,1,-1,2,0,-1,-1,1,0,0,-1,-3,1,-2,-1,0,0,0,0,0,-1,-2,-2,1,0,1,0,-1,-1,1,0,1,0,1,0,-1,-1,1,3,1,1,-1,-2,-2,1,0,0,1,0,0,0,1,-1,-3,1,0,1,-2,2,0,0,0,1,1,0,0,-1,1,-2,-1,0,-1,-1,2,-2,-1,2,-1,1,2,0,2,1,-2,0,0,-1,-2,1,-1,2,-1,0,-2,0,0,-2,-2,0,-1};
			304: counter1_out = '{-1,0,-1,0,0,0,-1,-1,1,0,1,1,-1,-1,0,-1,2,0,0,0,-1,1,2,0,0,0,1,0,-1,0,0,0,1,2,0,1,-1,0,0,-1,1,0,1,0,1,2,2,2,0,1,-1,1,1,0,0,0,0,-3,0,-2,2,0,-1,-1,1,0,3,-1,0,0,0,0,-1,-1,-1,2,0,-2,0,0,-1,2,-1,-2,-1,-1,0,-1,0,-2,3,-1,0,1,1,1,0,0,1,-1};
			305: counter1_out = '{1,0,0,-1,0,1,0,1,1,3,-1,0,0,1,1,-1,2,2,1,2,-1,0,-1,-1,0,2,0,-2,3,0,0,1,1,0,-1,0,-2,2,0,-2,1,1,0,0,1,0,0,2,0,-1,1,0,0,-2,1,0,1,-1,0,0,0,0,1,3,0,1,-1,-1,0,-1,0,0,2,-1,-1,-1,3,-1,1,0,-1,1,1,3,2,-1,0,0,0,1,-1,1,2,-2,2,0,-1,-1,-2,0};
			306: counter1_out = '{-1,-1,1,1,-2,-1,-1,0,0,2,0,0,1,0,0,-1,2,1,1,3,0,1,0,1,2,-1,-1,-1,1,-3,-1,0,1,-1,0,1,-1,1,1,0,1,0,0,1,1,-1,1,1,1,0,-1,0,1,-2,-1,1,1,-1,0,0,0,0,1,-1,-2,0,0,-1,1,1,1,2,0,0,0,-1,0,-1,-2,0,-1,0,-1,2,0,2,-1,0,1,1,-1,0,-1,1,-1,0,1,0,-2,-1};
			307: counter1_out = '{-1,-1,0,0,1,-1,-1,0,-2,-1,-1,0,-1,2,0,-2,1,-1,0,1,-2,0,2,1,1,1,1,0,0,0,1,1,0,0,-2,1,0,0,0,0,0,1,1,0,-1,2,1,1,-1,0,1,1,-1,-1,1,-1,0,-1,-2,-1,0,0,0,1,0,-1,0,-2,2,1,1,1,0,0,-1,0,1,0,2,0,-2,0,0,0,0,1,0,-2,2,1,3,0,0,-1,0,-1,-1,0,-1,1};
			308: counter1_out = '{1,0,0,0,-2,0,0,1,1,2,1,0,1,2,-1,-1,0,-2,0,2,0,1,0,0,0,1,0,0,0,0,-1,-1,1,0,0,0,1,-1,-2,-1,-1,0,2,1,0,0,-1,1,0,2,1,-3,0,-2,0,-1,1,0,1,-1,0,-1,-2,0,3,0,0,-1,0,0,-1,1,0,1,1,-2,1,1,1,0,0,0,-1,0,-1,0,-1,-2,1,-1,0,1,-1,1,-1,0,1,-1,1,1};
			309: counter1_out = '{0,1,2,1,0,-1,2,1,-1,-1,1,2,0,0,-1,0,-1,2,1,1,0,0,-1,-3,-1,1,0,-3,1,0,1,1,0,1,0,1,1,-1,0,-1,0,1,2,0,-1,3,0,0,-1,-1,-2,0,-1,0,0,-1,1,0,0,-2,-1,-2,0,0,0,0,1,1,1,0,0,1,2,0,-1,1,-1,-1,1,1,-1,-1,2,0,0,2,0,0,0,0,1,-1,-2,1,3,1,-1,-1,-1,1};
			310: counter1_out = '{-1,2,1,1,0,-2,0,1,0,0,-2,1,0,-1,-2,1,0,0,1,0,-1,0,0,0,0,-1,1,1,0,2,2,0,-1,-1,0,-1,0,0,1,-1,-1,0,0,1,0,1,1,-2,1,-3,0,2,-2,-1,-1,-2,0,0,1,0,1,1,1,-1,1,0,1,3,0,0,1,0,-1,-1,1,1,0,0,2,1,1,-1,-1,0,-2,0,0,-1,-1,1,-2,-1,-1,0,1,-1,0,1,0,0};
			311: counter1_out = '{-1,0,-1,0,1,-1,-1,0,-1,0,-2,0,1,-2,2,1,0,-1,-2,0,1,0,0,2,1,2,1,-1,0,-1,1,2,1,1,-1,-2,-1,-2,0,-1,2,0,2,1,0,1,-1,1,0,2,1,0,2,0,1,0,0,0,-1,0,0,0,1,0,-1,-1,-1,-1,2,-3,-1,0,-2,0,-1,-1,0,-1,-1,0,2,0,-3,1,-2,-1,-1,0,1,0,0,3,-1,0,1,0,1,0,0,0};
			312: counter1_out = '{-1,1,0,-1,0,0,-1,-1,0,0,0,1,-1,-1,2,0,2,0,0,1,1,1,0,0,1,0,-1,1,-1,0,-1,-2,1,0,0,-1,0,0,1,3,1,0,-1,-1,0,0,2,1,0,1,0,1,-1,-1,2,0,-2,-2,0,1,0,1,1,0,0,2,1,1,1,1,1,0,-1,0,0,0,-1,2,-1,1,0,0,1,1,-1,1,-1,-1,0,1,1,0,0,-1,-1,-1,0,1,0,0};
			313: counter1_out = '{-1,0,0,0,-1,1,1,0,-1,0,0,-1,0,-2,-3,-1,0,-1,-1,1,-2,1,-2,-1,-1,1,-1,0,-1,0,0,-1,1,1,1,0,0,-2,0,-1,-1,0,-2,-1,-2,0,-1,2,0,0,-1,0,0,-1,0,0,-1,1,-1,1,-2,0,0,0,3,-2,1,0,0,0,-2,0,1,2,-2,0,1,1,1,0,-1,1,-2,-3,2,-1,2,-1,2,0,0,0,-1,-2,0,0,-1,-1,0,2};
			314: counter1_out = '{2,-1,1,0,1,0,0,-1,0,-1,0,-2,0,-1,-1,0,2,0,-2,1,-1,-1,-1,1,2,-2,-2,-1,0,-1,1,-2,0,-1,-1,0,1,0,-1,-1,0,1,0,0,1,0,0,-1,1,0,0,0,0,1,-1,0,0,0,-1,1,1,0,-2,0,1,0,-1,0,0,-2,1,1,-2,0,-1,1,0,1,0,0,1,1,0,0,1,0,0,-1,2,1,1,-2,0,-1,0,-1,-1,0,0,0};
			315: counter1_out = '{-1,-1,1,-2,0,1,2,2,0,-2,-1,0,1,0,1,-1,0,-2,-1,0,1,1,-2,0,-1,0,1,-1,0,0,-1,0,-2,0,0,-2,-2,2,1,-1,0,0,-1,0,-1,0,0,1,-3,-1,-1,1,0,0,-1,1,1,1,1,2,1,1,0,0,-2,1,0,0,0,1,2,0,1,1,-1,1,1,-2,-1,1,0,1,-1,0,0,1,-3,-1,1,-1,0,0,-1,0,-2,0,-2,1,-1,-1};
			316: counter1_out = '{1,1,0,-2,1,0,0,1,1,-2,2,-1,0,0,-1,-2,0,0,-1,1,0,0,-3,1,-2,-1,0,1,1,1,1,-1,-2,0,-1,2,0,1,1,0,0,-1,0,0,-1,-1,1,-2,-1,-1,0,0,0,0,-1,0,1,-1,1,3,0,0,1,-1,-1,0,0,1,0,-2,2,0,-3,0,-1,0,0,-1,-1,1,0,0,1,2,0,-1,1,-1,2,-2,2,1,2,1,-1,0,-2,-1,1,1};
			317: counter1_out = '{-1,-1,-1,-1,1,-1,0,1,0,0,-3,0,0,2,2,-1,3,1,1,1,-2,2,-3,-1,-2,1,-1,0,0,0,0,1,-1,2,-1,-1,-1,0,3,-2,1,1,-2,-1,-1,1,2,1,-2,0,-1,0,0,-1,-3,-1,0,1,2,2,1,1,0,-1,0,-2,-1,0,2,0,1,1,1,0,0,2,0,-1,-1,1,-2,0,1,2,1,0,-1,0,1,0,0,0,0,1,3,0,-2,-1,-1,1};
			318: counter1_out = '{0,-1,2,2,-2,-2,-2,1,-1,-2,-2,0,1,0,1,1,2,4,-1,1,-2,1,-3,2,0,0,-1,-1,1,0,-2,1,-1,0,-1,0,0,0,2,-1,1,2,0,0,0,1,0,1,0,0,-1,0,-2,2,0,0,-1,0,1,1,-1,0,1,-1,-1,-1,0,0,0,-1,1,0,-1,1,-2,0,2,0,1,-1,-2,1,0,0,1,0,-3,0,1,1,0,-1,0,0,-1,2,-1,-1,0,0};
			319: counter1_out = '{-1,-2,0,2,-1,-2,-1,1,1,1,0,0,0,-1,2,0,-1,1,-1,0,-1,1,-4,-1,-2,0,-1,-1,1,-1,0,1,-1,1,-1,2,-2,0,0,-1,-1,0,-1,-1,0,0,-2,-1,0,-1,-2,1,2,1,0,1,-1,2,-1,2,0,1,0,-1,-1,1,-1,0,1,-1,1,0,-2,2,-1,2,2,0,1,1,1,1,1,1,2,1,0,0,1,0,0,0,-2,0,1,0,-1,-2,-2,0};
			320: counter1_out = '{-1,-1,1,1,0,-1,0,0,-1,0,-1,-2,0,-1,-1,1,1,1,0,1,-3,0,-2,1,-1,0,0,1,2,0,0,1,-1,0,0,0,-2,-1,-1,1,1,-2,-1,-1,-1,-1,-1,0,1,1,-1,1,0,-1,-2,-2,-1,1,1,0,2,2,1,1,0,0,-1,-2,0,1,1,1,-1,-1,-1,1,2,1,1,-1,-1,1,1,0,-1,1,-4,0,-1,1,0,1,0,0,1,0,-3,-1,1,-1};
			321: counter1_out = '{-1,1,1,2,0,-2,0,0,-1,1,-2,-2,-1,-3,-1,1,0,-2,1,1,-1,0,-2,0,-2,0,1,-1,2,-1,2,1,-1,1,2,1,-3,0,-1,1,-1,-1,-2,0,-2,1,-1,1,2,-1,0,0,0,-1,2,-3,0,0,0,1,0,1,-1,0,-2,-2,0,0,0,0,1,-1,0,-1,0,1,-1,0,-1,-1,0,1,2,0,2,0,-1,1,0,0,0,0,1,0,1,1,-4,-1,0,-1};
			322: counter1_out = '{1,2,2,0,2,-3,0,-1,1,0,0,-2,0,-1,0,1,-2,-1,1,0,0,0,0,-2,0,0,0,-1,0,2,-1,1,1,-2,2,-1,0,-1,-1,1,2,-2,0,-1,-1,2,-2,0,1,0,1,-1,1,1,1,-1,2,-2,1,0,0,-2,0,-1,0,0,0,1,2,1,1,0,1,-1,-1,2,1,-1,1,1,0,1,2,0,0,-1,-3,1,3,1,0,1,0,-2,-2,0,0,-1,-1,2};
			323: counter1_out = '{1,2,1,2,1,1,1,1,1,1,-1,1,0,-1,0,1,0,-2,0,0,1,-2,0,0,0,-1,-1,-2,0,-2,0,0,0,0,1,-1,2,0,-2,2,2,-1,1,-1,-2,-1,1,2,0,-1,1,-3,1,1,1,0,1,-2,1,1,-1,0,0,0,-1,-2,-2,1,1,1,0,0,0,1,0,-1,2,2,0,1,0,1,3,0,-2,0,1,1,1,-1,-2,-1,0,-1,-3,2,1,0,0,2};
			324: counter1_out = '{0,0,-1,0,1,-1,-3,0,0,1,0,-1,1,-1,1,-1,3,1,-1,-1,1,2,-1,0,-1,-2,-1,0,1,-2,-1,-1,1,0,-1,-1,1,-3,-1,2,1,-1,0,-1,0,0,0,0,0,1,1,-3,1,0,1,1,0,1,0,0,2,0,0,1,2,-1,1,0,1,-2,0,1,-1,-1,-1,-1,0,2,0,-1,-2,1,-1,1,1,1,-1,0,-2,-2,-2,0,1,-1,-2,1,-2,0,2,2};
			325: counter1_out = '{1,0,-1,1,0,-1,2,-1,-1,-1,-2,-1,0,-1,0,1,0,2,1,1,-1,1,1,0,0,-1,-1,0,1,-1,0,-1,0,1,0,0,1,0,1,0,0,0,0,1,-1,0,-2,1,-1,0,0,-1,0,0,-1,1,-1,-1,2,0,1,-1,-1,-1,-1,0,1,3,0,-1,0,1,0,-1,-2,1,2,0,-2,0,1,-1,-1,0,2,1,0,-1,1,-2,0,-1,0,0,2,4,0,-1,0,1};
			326: counter1_out = '{0,0,-1,-1,0,0,2,1,-1,-2,1,-4,0,-2,3,-1,0,1,0,0,1,1,1,0,0,-2,0,1,1,0,1,-2,-2,0,-1,1,0,-4,-1,0,1,1,1,-1,-1,2,1,1,-2,1,1,2,0,0,-1,0,0,-1,1,-1,-1,1,0,0,-1,0,1,1,2,1,1,3,-1,1,-1,-1,-1,-1,0,1,0,1,-2,0,0,3,0,0,-1,0,-2,-1,0,0,1,2,1,2,1,1};
			327: counter1_out = '{-1,1,0,-1,1,0,2,-1,0,-1,-1,0,1,0,0,-1,0,-1,0,0,-1,-1,3,-1,-1,-2,3,-2,-1,0,1,-1,1,0,0,-1,2,-3,-1,3,0,-2,1,-1,-1,0,0,0,-2,0,0,1,3,-1,2,0,-1,1,1,-1,1,-1,-2,1,-1,0,2,-1,0,-2,1,1,1,1,1,2,-1,-1,1,-2,0,-1,0,0,0,0,0,-1,0,-2,-1,2,-1,1,1,2,1,-1,0,1};
			328: counter1_out = '{-1,0,-2,-1,1,0,1,0,1,-2,0,-3,1,0,0,1,-1,-2,0,2,-1,2,0,0,1,-3,1,0,1,2,-1,-2,1,-1,0,2,3,-2,-1,0,-2,-2,0,-2,1,1,2,1,-2,-2,2,2,1,0,0,-2,0,-1,1,0,1,1,-1,1,-1,1,2,1,0,-1,1,1,1,-1,1,-1,0,1,-1,-1,0,0,-2,0,0,1,0,0,2,-3,-1,2,-2,1,1,1,1,-1,0,2};
			329: counter1_out = '{1,1,1,1,1,1,-1,3,0,0,0,0,0,1,0,1,-1,1,2,2,-1,1,-1,-1,0,-2,1,0,-2,0,2,0,0,1,-1,-1,-1,-1,0,-1,1,1,1,0,0,3,1,1,1,1,3,1,0,-1,0,0,0,-1,-1,0,0,-2,-2,0,1,1,2,-1,0,0,0,0,0,0,0,0,0,-2,-2,2,-2,-1,0,0,-1,0,-1,0,2,0,0,1,0,0,-1,1,-2,0,-2,-1};
			330: counter1_out = '{0,1,1,-2,-1,1,0,0,1,2,-1,-1,0,2,1,-2,-1,-2,0,0,-2,1,0,0,0,-1,-1,0,0,0,1,2,-2,0,0,-1,-1,-1,1,-3,-2,1,0,-1,0,1,-1,2,-2,-1,0,-1,-1,-2,-1,-4,1,-1,1,0,0,1,-1,-1,-1,-1,0,1,0,-1,0,1,2,0,0,0,-2,0,0,-1,1,-1,0,1,-2,0,-1,2,1,-1,1,-1,1,1,0,3,1,1,1,1};
			331: counter1_out = '{1,-2,2,-1,0,-2,2,1,0,0,-1,0,1,0,-1,0,1,-1,0,0,0,0,-2,0,-3,1,1,1,-1,0,2,0,0,1,0,-1,-2,0,0,-2,0,0,0,-3,0,-1,0,0,-2,-1,-1,0,0,-1,0,-1,0,-1,-1,0,0,-1,1,-3,-1,-1,-2,1,1,1,-1,-1,-2,1,0,1,-1,0,-1,-1,1,-1,1,-1,0,-1,-3,0,0,0,1,0,0,0,2,2,0,1,0,1};
			332: counter1_out = '{0,0,0,-1,-1,-1,0,1,2,-1,-1,0,1,-2,-2,-2,1,-2,2,1,-1,0,0,0,0,1,0,0,1,0,-1,1,0,-1,0,2,-1,0,1,-1,1,1,2,-1,1,0,-2,1,0,-1,-2,0,0,-2,-2,-2,1,0,2,0,0,0,0,1,-1,1,-1,0,0,1,1,0,0,0,1,-1,2,1,-1,1,-2,0,0,-1,-2,0,-1,-1,1,-1,1,-1,1,0,1,1,0,-2,0,2};
			333: counter1_out = '{2,0,-1,0,-1,0,-1,0,2,0,-1,1,1,1,0,-1,0,2,0,-2,-1,1,1,0,0,1,1,-1,-2,1,1,2,0,0,0,-1,1,0,-1,-1,2,1,-1,1,1,-3,1,1,0,2,2,2,-2,0,1,0,2,-1,1,1,-3,0,-2,0,1,-1,0,-1,-1,-1,0,-1,-3,-1,2,1,2,0,1,0,2,0,1,-1,1,0,0,-3,0,-1,-1,-1,0,-1,3,-1,0,1,1,-2};
			334: counter1_out = '{1,0,-1,1,-1,0,-1,-2,1,0,0,0,-1,0,2,3,0,1,-1,0,1,2,1,-2,1,1,0,-1,0,0,0,0,1,0,2,0,0,-1,0,0,-1,0,-1,0,-2,-1,-2,-1,-1,0,0,0,1,1,1,1,0,-1,1,2,-1,0,0,0,1,-1,0,-1,0,-1,0,-1,-1,0,0,1,1,-1,0,0,0,0,1,-1,-2,0,-1,-1,0,1,-1,0,-1,0,0,2,1,-1,0,-1};
			335: counter1_out = '{1,1,1,0,0,-1,-1,-1,0,-1,1,0,1,0,-1,0,1,-1,-1,0,0,0,1,-2,-1,2,0,0,1,0,-1,0,-1,0,0,1,-1,-2,0,3,2,0,1,0,0,1,0,1,1,0,-1,0,2,0,0,0,0,1,-1,2,0,1,2,1,1,-1,1,0,-1,1,-2,2,0,1,2,0,0,1,-1,-1,-1,0,-3,2,1,-1,2,0,-1,1,2,0,0,1,0,0,1,1,1,-1};
			336: counter1_out = '{2,-1,1,0,-2,0,-2,0,0,-1,1,1,1,-1,-1,1,1,0,0,0,0,0,0,1,0,-1,-1,0,-1,0,-2,1,0,1,1,1,-1,2,0,2,1,1,-1,-1,1,2,0,1,1,1,1,-1,-2,1,0,1,0,1,0,-1,0,0,-1,0,1,-1,0,-1,2,0,0,1,-2,-1,-1,0,0,1,0,0,0,-3,0,0,0,0,1,0,1,1,0,-1,-1,1,1,1,-1,2,0,1};
			337: counter1_out = '{-1,0,0,2,-1,0,-1,-1,0,-2,0,0,-1,-1,0,1,-1,0,0,2,1,-1,0,0,0,-1,0,0,0,2,1,0,1,0,-1,1,1,0,-1,0,0,0,1,0,3,0,-1,0,-1,2,0,0,2,0,2,1,1,1,0,-2,-2,2,-2,-1,1,1,-1,0,-1,-1,1,1,1,0,0,0,-1,0,-1,-1,0,-1,-1,2,1,1,-2,0,1,0,0,0,-2,0,0,0,-1,-1,0,-2};
			338: counter1_out = '{0,1,0,0,0,0,0,1,0,-1,-1,-2,1,1,0,0,1,0,0,-1,0,0,1,3,1,1,0,0,-1,0,0,0,1,2,-2,0,-1,1,0,0,0,-1,0,1,0,0,-1,2,0,0,-3,1,0,0,0,0,1,1,1,0,-2,-1,-1,-1,1,0,-2,0,0,-2,0,-1,1,0,0,-1,1,-3,0,1,0,1,0,0,-1,-2,2,1,-1,1,1,0,-1,-1,2,-1,0,-2,-1,-1};
			339: counter1_out = '{1,0,3,-1,-1,-2,0,0,-2,0,1,-1,1,0,-1,2,0,1,1,-1,0,1,-1,0,0,2,1,2,-1,1,1,0,0,0,-2,-1,-1,1,0,1,-1,-1,0,0,-2,-2,0,0,0,0,2,0,0,0,0,2,-1,0,1,1,-1,0,1,-1,0,-1,-1,1,2,0,0,-1,-1,0,1,1,1,-1,1,0,1,0,0,2,0,1,-1,0,2,0,1,0,0,1,2,1,0,2,-1,0};
			340: counter1_out = '{0,-2,1,1,1,0,1,1,0,0,-2,-1,1,0,-1,0,0,0,-1,0,-1,2,-1,0,1,-1,0,0,0,-1,1,0,1,1,-2,0,-1,1,1,2,0,1,1,-2,0,-2,1,1,-1,-1,0,-1,0,-2,1,-1,0,0,1,-2,-1,-1,1,0,2,-2,0,1,1,0,-1,3,1,0,0,-1,0,-1,-1,1,0,-1,-2,-1,0,2,-1,0,-1,1,0,1,-1,-1,1,1,-3,0,1,0};
			341: counter1_out = '{-1,-1,0,0,1,-2,-1,0,1,1,0,1,1,2,0,-3,0,-2,-1,1,-1,-1,-2,0,-1,0,1,1,-1,0,-1,-1,-2,-1,2,-1,-2,-1,3,-1,1,0,0,1,1,1,-1,1,-2,0,1,2,-2,-1,0,0,-1,0,0,0,2,2,1,-1,-1,1,-1,0,2,-1,-2,1,0,-1,-1,-1,1,-1,1,1,0,1,0,0,-1,0,-1,-1,0,-1,1,0,-1,0,-1,0,-3,0,-1,2};
			342: counter1_out = '{0,1,0,0,1,0,-2,0,-1,-1,1,1,0,0,-1,0,1,1,0,2,-1,0,-3,0,0,0,1,-1,0,-1,0,-1,0,1,-1,0,0,1,0,1,-1,0,0,-2,0,0,-2,1,-1,0,-2,1,-1,0,0,1,0,-1,-1,0,1,0,0,-1,-1,-1,2,-1,-1,1,-2,1,-2,0,-1,0,1,-1,0,-1,-1,1,-1,0,0,-2,-1,0,0,-1,2,0,0,-1,-1,-1,-1,0,0,-1};
			343: counter1_out = '{-1,-1,0,-2,0,-1,0,0,0,-1,1,4,1,1,1,0,2,0,-1,1,1,-1,-3,0,-1,1,0,1,0,1,0,0,-3,-1,0,-2,0,-1,1,0,1,0,2,2,1,0,2,0,-1,-1,1,1,0,-2,0,0,2,0,2,0,-1,-1,1,0,1,-1,0,0,-1,1,1,-1,1,-1,1,0,-1,3,1,2,2,-1,1,1,0,1,-2,1,-1,0,0,0,0,-1,0,0,-1,0,0,1};
			344: counter1_out = '{-1,-1,-1,1,0,0,0,2,-2,0,-2,0,1,1,1,0,0,1,-1,0,0,1,-3,0,-2,-1,-1,-1,1,-3,0,0,1,0,-2,-1,0,0,3,1,0,1,-1,-1,1,-1,0,-1,-1,1,-1,0,1,0,0,0,-2,1,1,-1,0,0,-1,0,1,1,1,0,-1,0,1,0,-1,0,0,1,0,0,0,-1,-2,1,-2,0,1,0,-1,0,0,-2,-1,-2,1,0,1,0,0,-1,0,0};
			345: counter1_out = '{0,0,0,0,0,0,-1,1,0,-1,1,1,2,0,-1,1,2,2,0,1,-1,-1,-5,-2,-2,0,0,1,0,0,0,0,0,0,-1,0,0,0,1,0,0,0,-2,1,1,1,0,-1,0,0,0,1,-2,1,-2,-1,-1,0,1,0,1,1,0,-1,-2,-1,1,1,-1,-1,-2,-1,1,-1,1,2,1,1,-1,0,0,2,-3,-1,0,3,-3,-2,2,-1,0,0,-1,-2,0,1,0,-1,-1,0};
			346: counter1_out = '{0,0,2,0,0,1,0,1,-1,1,2,0,2,-1,1,0,-1,2,0,0,1,1,0,0,-1,-1,0,1,1,1,-1,0,1,-1,-1,0,1,0,0,0,1,2,0,0,0,-1,-2,1,2,0,-1,1,-1,-1,0,-1,1,1,1,-2,0,2,-1,0,-2,0,-1,0,-2,1,2,0,2,1,1,2,0,2,-1,0,0,0,0,0,0,0,0,0,-1,2,0,-1,0,1,0,-1,0,-2,1,0};
			347: counter1_out = '{1,0,1,2,-1,0,-3,0,0,1,-1,0,2,0,0,1,-1,1,1,0,0,2,0,1,-1,1,1,2,2,-1,1,1,-1,0,-1,1,0,0,-2,0,-2,4,-1,1,-1,0,-2,0,-1,0,-1,2,-1,-1,-1,1,-1,1,-1,-1,2,1,0,0,-1,-2,0,1,-1,1,0,2,-1,1,0,0,-1,1,-1,1,-1,-1,-2,-1,1,-1,-4,1,0,0,1,0,1,1,1,2,-1,1,0,0};
			348: counter1_out = '{-1,-1,-1,1,-1,-2,2,-2,0,1,0,-2,2,0,0,1,-1,-2,-2,0,-1,0,1,0,-1,0,-1,0,0,-1,2,-2,1,1,-2,2,0,0,-2,-1,2,1,0,0,-1,-2,-2,1,0,0,-1,-2,-1,1,-1,0,0,0,2,-1,0,3,1,0,-1,-1,-1,0,0,-1,-1,1,0,0,2,3,1,0,2,-1,0,0,-1,-2,1,-1,-2,1,-2,-2,2,1,-2,0,1,0,-2,1,1,-1};
			349: counter1_out = '{2,-1,0,0,0,-1,1,-2,-2,-1,0,-2,0,0,1,0,0,0,1,1,0,0,0,-2,-1,2,0,0,2,1,2,1,0,3,1,1,-4,3,-1,0,1,-1,-1,0,-1,-1,-2,0,1,-1,0,0,2,0,0,0,-1,-1,0,-1,-1,0,1,-1,-1,-1,1,1,0,1,0,3,0,-2,1,2,1,1,0,0,-1,0,-1,-1,-1,0,-2,1,2,1,2,1,-1,0,-1,2,2,-2,0,-1};
			350: counter1_out = '{4,0,0,0,1,1,1,-1,0,1,-1,-1,1,-1,0,0,-2,0,0,0,-2,-3,0,0,1,0,-1,-1,0,0,1,1,-1,1,2,0,1,0,-1,1,0,-2,1,-1,-1,-1,0,0,2,0,2,0,2,1,1,-1,1,-1,-1,0,0,1,0,0,-2,-4,-1,0,-1,1,1,0,0,0,0,1,3,1,-1,0,-1,-2,0,-2,2,-1,-1,0,2,1,0,0,-1,-2,-3,1,1,1,0,0};
			351: counter1_out = '{1,1,3,0,-1,0,-1,-2,0,-1,0,-2,-1,-1,-1,0,-1,-1,1,0,-1,1,-2,-1,0,0,0,-2,0,-2,0,1,1,2,2,0,2,-1,-1,0,0,0,1,0,-2,-1,0,1,1,-1,1,-1,0,1,2,1,1,0,0,0,0,0,-1,0,0,-2,1,2,-1,1,1,1,0,0,-1,1,2,2,-2,0,1,-1,0,1,0,-1,0,0,2,-1,-1,2,-1,0,0,0,2,1,1,1};
			352: counter1_out = '{0,1,0,1,0,1,-2,0,-2,0,-1,0,0,0,0,-2,0,0,-2,2,1,-1,1,-1,0,-1,1,-1,-1,-1,1,0,0,-1,0,0,2,-2,0,-1,0,1,0,1,-3,0,1,1,0,-1,1,-2,-2,-1,-1,-1,1,0,-1,0,1,1,0,0,-3,-1,0,0,-3,0,-1,0,-1,-2,-1,2,0,-1,-2,-1,1,1,0,0,1,2,-2,0,1,0,-2,1,0,1,0,2,0,0,-2,0};
			353: counter1_out = '{-2,0,-1,1,0,1,1,-2,-1,0,-1,0,-1,-2,1,1,-1,1,-1,0,-1,0,-1,1,0,1,-2,-1,-1,-1,-1,1,-1,0,-1,2,3,-3,0,-1,-1,-1,-1,0,0,0,-1,-1,-1,-1,1,-2,-1,-1,-1,0,1,1,2,1,1,-1,-1,0,0,0,2,1,-1,0,-1,0,-1,0,-1,1,-1,-2,-1,-1,0,0,0,-1,1,0,-2,0,0,0,-2,2,0,-3,1,1,0,0,-2,-1};
			354: counter1_out = '{-2,-1,0,2,1,0,0,-1,-1,1,1,0,-1,-1,-1,-2,0,-1,-1,0,-1,1,0,0,0,-1,-2,-1,1,-1,-1,-2,-1,0,0,0,0,-3,-1,-1,1,-2,0,-4,-2,1,1,0,-2,1,0,0,1,0,-1,-1,-1,1,1,-2,0,-2,0,0,1,-2,0,2,0,-2,1,0,-2,0,-2,-1,1,1,-1,-1,1,0,-1,-1,0,0,0,1,1,-1,0,1,0,0,1,1,0,-2,1,0};
			355: counter1_out = '{0,-1,0,0,0,1,1,0,1,1,-1,-1,0,0,2,1,-1,1,-2,2,0,1,0,1,-1,0,1,0,-1,0,1,-2,0,-1,1,-3,1,-2,0,-1,0,2,-1,1,0,1,1,-1,-1,0,0,1,-1,0,1,0,0,2,1,-2,0,0,-1,1,1,0,1,0,0,1,2,0,1,-1,-2,1,-1,-1,1,-2,1,2,-1,-1,1,0,-1,-2,1,-1,-1,1,-3,-2,1,2,3,1,-1,0};
			356: counter1_out = '{0,-1,-2,2,0,0,0,-1,-1,-1,0,-1,-1,1,1,1,-1,1,4,1,0,0,0,0,0,0,0,0,0,-1,-1,0,0,-1,-1,-1,0,-3,-1,-2,0,0,0,0,1,1,-2,0,0,-1,0,0,2,-1,0,-2,0,1,1,0,1,-1,1,-1,0,1,1,1,0,-1,-1,0,0,0,-1,0,1,1,1,-1,0,1,0,1,-1,0,-1,2,0,-1,-1,1,-1,0,0,0,0,0,0,0};
			357: counter1_out = '{0,-1,-1,-1,-2,1,1,0,0,0,1,0,0,0,0,-1,2,1,-1,1,0,0,0,-1,0,0,1,2,1,0,1,0,0,0,-1,1,0,-3,0,-2,0,-1,1,0,0,1,-1,1,-1,-1,0,1,-1,-1,-2,-1,1,1,2,-1,0,1,0,-1,0,2,1,0,1,1,1,-1,1,0,2,0,-1,-1,-1,-1,0,0,1,0,1,0,-3,1,-1,0,-1,0,1,1,1,1,0,-1,1,0};
			358: counter1_out = '{1,-1,-1,2,-2,2,0,0,0,-1,1,-1,1,0,0,-1,-2,2,0,1,1,0,0,1,2,-1,-1,-1,0,2,-1,0,-1,-2,1,0,0,-2,-1,-2,-2,-1,1,-1,0,2,3,1,-1,-1,0,3,2,-2,0,-1,2,0,2,0,0,1,1,0,-1,1,2,0,2,-1,0,-1,0,2,0,-1,0,2,0,0,0,0,-1,-1,2,0,-2,0,-1,0,-1,-1,0,-3,-1,0,-2,0,-1,1};
			359: counter1_out = '{1,0,-1,1,1,1,1,-2,-1,1,0,0,0,0,1,-2,-2,0,0,0,1,-1,1,0,-1,1,0,1,2,0,0,0,-1,0,-2,0,0,-3,0,0,-1,-1,2,-1,0,-1,0,3,0,-2,-1,3,-1,1,-2,0,2,2,0,-1,-1,-1,1,-1,0,1,0,2,0,1,1,0,-1,1,0,0,0,0,1,-1,1,2,0,0,0,0,-2,1,1,-1,0,0,0,-2,-2,0,0,-1,-1,2};
			360: counter1_out = '{1,-2,-1,0,1,1,-1,-1,1,-2,1,-1,-1,-1,-1,-1,1,-1,1,2,0,0,0,1,-1,0,0,1,0,0,-1,0,2,1,0,-1,-3,-4,0,-1,-3,1,1,-1,0,-2,1,0,1,-1,0,-2,0,1,0,0,-1,0,1,-1,-1,1,-1,-2,-2,1,-1,0,1,-1,0,-1,0,-1,1,1,-1,-1,0,0,-2,-1,1,0,0,0,-1,0,-1,1,1,1,0,0,-1,3,-3,0,-2,0};
			361: counter1_out = '{-2,-2,-1,-1,1,0,0,-2,0,-1,0,-1,0,2,0,1,0,1,1,-2,-1,-1,1,-2,0,1,1,0,1,-1,1,-1,2,0,2,0,-1,-1,1,-1,-2,1,-1,1,0,0,1,0,1,-1,1,1,0,-2,0,0,0,0,1,0,0,-1,-1,-1,0,0,1,1,0,-1,-1,0,2,0,-2,0,0,0,-1,0,1,0,0,0,-2,-1,-1,0,0,0,0,0,0,1,1,0,-1,0,-2,0};
			362: counter1_out = '{-1,2,0,0,0,0,1,0,0,0,1,-1,-1,0,-2,-1,-1,1,2,0,0,-1,0,-1,0,-2,1,1,0,0,0,1,1,0,0,0,1,1,1,-2,-1,-2,0,-1,3,0,-2,-1,0,-1,0,0,0,0,2,-1,2,0,-2,2,0,1,-1,0,0,1,0,1,0,-1,0,-1,-1,1,-2,0,0,-1,-1,0,1,-1,0,1,1,0,0,1,0,2,0,-1,1,0,1,2,-1,1,-1,2};
			363: counter1_out = '{0,0,1,0,-1,-1,-2,0,1,-1,0,-1,0,1,-1,1,-1,0,0,1,-1,1,0,1,1,-1,0,-1,1,-1,-1,1,0,0,-1,0,1,-1,1,0,-2,1,-2,0,-1,-1,1,1,0,0,1,0,-1,-1,0,0,1,0,1,-1,1,-1,-2,0,-2,-1,0,0,1,2,1,-1,1,0,2,1,0,0,1,1,-1,0,-1,0,-1,0,-1,-1,0,1,0,1,0,0,1,0,1,0,0,1};
			364: counter1_out = '{-1,-1,0,-1,-1,0,0,-1,0,-1,-1,2,-1,0,0,0,0,1,0,0,0,1,0,-1,0,-2,2,-1,1,1,1,0,1,-1,0,0,-1,0,0,1,0,0,0,0,1,1,1,0,1,0,-2,0,1,1,0,1,1,-2,0,0,0,0,1,-1,1,0,0,1,0,0,-1,0,0,-2,1,0,-1,0,-1,2,-1,0,0,0,-1,1,1,1,-3,0,0,0,-2,0,0,-1,0,0,0,0};
			365: counter1_out = '{1,0,0,-1,0,1,0,1,0,0,0,1,1,0,-2,0,0,-1,-2,-1,-2,1,-1,-1,0,0,-1,1,0,-1,0,1,0,1,1,0,0,-1,1,0,-1,1,-1,1,1,0,1,1,0,-1,1,0,0,1,-2,0,-1,-1,0,-1,0,1,-1,2,0,0,0,0,0,0,0,-1,0,0,0,0,0,-1,0,2,0,0,1,1,1,-1,0,-1,-1,2,0,-1,-1,-3,-1,0,-1,1,-1,-1};
			366: counter1_out = '{0,1,-1,1,0,1,0,-1,1,-1,1,0,3,-1,1,1,0,-1,0,-1,0,-1,1,-1,1,-1,-1,0,1,1,-2,0,-1,0,2,0,1,-1,1,0,-1,0,-1,-2,-1,1,1,1,-2,2,0,0,1,0,1,1,0,-1,0,-1,-1,0,1,0,-2,-1,-1,-1,0,1,0,-1,-1,1,0,-2,0,0,1,0,0,2,0,0,0,0,-1,1,0,-1,-1,1,0,0,-1,0,0,0,1,0};
			367: counter1_out = '{0,-1,1,0,1,0,0,0,0,1,-1,0,1,1,1,-1,1,0,1,-1,1,-1,-1,0,0,-1,0,-1,0,-1,0,1,0,1,1,1,2,1,1,0,-1,0,-2,0,0,-2,1,-1,0,0,2,0,1,1,0,0,-1,-3,0,-1,-1,-1,0,-1,1,-1,-1,2,0,3,0,-1,0,1,-1,0,1,1,2,0,0,0,-1,1,1,1,1,0,-1,0,-2,1,-1,0,0,-2,0,-2,0,1};
			368: counter1_out = '{-1,1,0,-1,0,-1,1,-1,1,0,1,-1,-2,1,-1,-1,2,2,1,-1,1,2,-1,0,-2,0,0,2,1,-1,0,-1,0,1,1,1,0,-1,1,-1,-1,1,0,1,0,1,0,1,0,0,-1,3,0,0,1,-1,1,2,1,1,1,0,0,0,1,0,-1,0,1,-2,1,-1,0,1,-1,1,-1,-2,0,-2,0,4,-1,0,0,0,-2,0,0,2,-1,1,0,-1,-1,0,0,1,-1,0};
			369: counter1_out = '{-1,-1,3,-3,0,0,1,-1,-1,-1,0,1,2,-2,-1,-1,1,0,1,0,-2,0,-3,0,-1,-2,0,0,1,-1,-1,-1,0,0,-1,-1,0,0,0,0,1,0,-1,-3,1,-1,2,0,-1,-1,-1,1,0,-1,-2,0,-1,-1,0,0,0,3,0,2,0,0,-1,1,1,-2,0,1,-2,0,-1,-1,-1,0,0,0,1,1,0,0,-1,2,0,-1,1,0,0,0,0,-1,2,1,-2,-2,-1,2};
			370: counter1_out = '{-1,-1,0,0,0,0,-1,-1,-1,2,-1,2,1,-1,-2,-1,1,0,-1,1,0,1,-1,1,-2,0,1,1,1,1,-1,0,-1,0,-2,0,1,-1,1,-1,0,2,1,-1,-1,0,1,-1,1,0,0,0,0,1,-2,1,0,1,0,0,1,2,1,0,-1,0,1,1,1,1,3,-1,0,1,-1,0,0,0,1,-1,0,0,-2,0,0,-1,-1,-1,-1,0,1,-2,0,1,-1,-1,1,0,1,0};
			371: counter1_out = '{1,0,-1,1,-1,-1,0,2,0,2,-2,-1,-1,0,-1,-1,2,1,-2,1,0,1,-2,-1,-1,-2,0,1,2,2,1,-1,0,0,-4,0,1,2,0,-1,1,0,1,1,0,2,-1,1,1,-1,1,0,-1,0,-1,0,0,1,1,0,0,-1,0,0,-2,-1,0,-1,0,0,-1,2,-1,1,0,0,0,0,-1,1,-2,1,-2,0,0,1,-3,1,0,1,-1,-1,1,1,-1,2,-1,-1,0,0};
			372: counter1_out = '{-2,-1,3,0,-1,0,-1,1,0,0,0,0,1,0,1,0,0,0,-2,2,1,-1,-2,-1,-2,0,1,0,1,1,-2,0,0,1,-1,2,-1,0,1,-1,-1,1,-2,-2,-1,0,0,1,-1,1,-1,0,0,-3,0,-1,1,0,1,-1,0,1,-1,3,-2,0,0,0,-1,2,0,0,1,0,1,1,-1,1,1,1,0,-2,-1,-1,0,0,-2,-2,0,-2,2,0,-1,1,-1,1,0,-1,0,-1};
			373: counter1_out = '{0,0,0,-2,0,-1,0,0,-1,3,1,2,1,-2,2,1,1,2,-1,2,1,1,3,0,-2,-1,1,1,2,-1,-3,1,-1,0,-2,2,0,0,4,-1,-1,1,1,0,-1,1,0,1,0,0,0,0,-2,1,-1,0,-1,-1,0,-1,0,0,0,0,-2,-1,0,-1,-2,-1,1,-1,1,1,1,3,1,-1,0,0,0,-2,-2,0,0,-1,-1,2,2,-2,1,0,1,0,1,0,-1,0,-2,0};
			374: counter1_out = '{-2,-1,2,0,2,-1,-1,-1,1,2,0,0,0,-1,1,1,0,0,-1,-1,0,1,1,-2,-2,-1,0,0,1,1,-1,1,0,0,-1,0,-2,1,2,-1,1,2,0,1,-1,-1,-2,0,-1,2,-1,-1,0,0,0,1,-2,2,1,-1,-1,1,-1,0,-1,-1,-1,0,0,-1,-1,0,0,0,0,1,1,0,0,0,0,0,-2,0,1,0,0,0,0,1,-1,-2,1,1,1,2,-1,-1,2,0};
			375: counter1_out = '{-2,0,0,2,0,0,0,-1,-2,2,0,-1,2,-1,2,1,-1,-1,-2,-1,-1,1,-1,0,-1,1,0,0,0,2,-1,0,-1,0,-2,1,0,-1,1,0,0,2,0,-2,-1,-1,-2,0,1,-1,0,1,1,-2,-2,0,-1,1,-1,1,0,0,1,-1,0,1,0,-1,-1,2,0,-1,-1,0,1,1,2,-1,1,-1,1,1,-3,-2,1,0,-1,0,1,1,0,1,0,1,0,1,-1,1,-1,1};
			376: counter1_out = '{1,-1,0,1,-1,0,1,-3,-1,0,0,0,2,-2,0,0,0,-2,1,0,-2,-1,0,1,1,0,0,2,1,0,2,1,1,3,-3,1,-1,1,0,0,1,3,0,1,0,-3,-2,-2,0,1,0,-2,-1,-2,0,-2,1,-1,1,-1,0,1,1,-1,0,-2,1,0,1,1,1,1,1,-1,0,0,0,-1,-1,1,0,-1,-3,-1,0,-2,-2,0,2,1,3,0,1,1,-1,0,-1,0,0,0};
			377: counter1_out = '{2,0,1,1,0,-2,2,-1,0,1,1,0,1,-1,0,2,1,0,1,1,-1,1,1,0,1,0,-1,0,0,-1,0,2,0,0,1,2,0,-1,0,1,1,0,-1,-1,-1,-1,0,1,2,-1,0,0,1,1,1,0,1,0,-3,0,-2,1,1,-1,1,-2,0,1,-1,2,-1,0,-2,-4,0,0,0,2,0,0,0,1,-1,3,0,0,1,1,1,1,1,0,1,1,-1,-1,-1,0,-1,-1};
			378: counter1_out = '{4,0,0,0,2,-1,0,0,0,0,1,0,-1,0,0,0,1,0,1,0,-1,0,0,-3,1,1,-1,1,1,-1,2,1,-1,0,0,3,2,-1,1,1,1,-2,1,-1,0,0,-1,-1,1,0,1,-1,0,0,0,0,0,0,-1,2,-1,-1,1,0,-1,-1,-1,0,-1,-1,-1,-1,1,0,-1,1,1,0,-1,0,1,0,-3,-1,2,-1,0,1,1,3,0,2,1,-3,-1,0,-2,0,0,1};
			379: counter1_out = '{2,1,2,0,0,1,-1,0,-1,-2,0,-1,-3,-1,0,0,2,-2,-1,0,-1,1,0,0,-1,0,0,1,0,-1,1,0,-2,2,2,0,0,-2,0,1,-1,0,0,0,-1,0,1,0,-1,-1,1,1,0,1,-2,0,0,2,1,-2,-1,2,0,2,0,0,-1,0,-2,-1,0,0,0,0,-2,1,0,0,1,0,-1,-2,-2,0,2,1,1,-1,1,-2,-2,1,0,-1,-2,0,-1,1,-1,1};
			380: counter1_out = '{0,-2,0,0,-1,-2,2,-2,1,1,0,0,-1,0,1,0,0,0,0,0,0,1,-1,0,-1,1,-3,-1,1,-2,0,0,-1,0,1,-1,1,0,0,0,0,0,0,1,1,-1,0,1,0,1,0,-2,2,1,0,0,1,1,1,0,0,-1,-2,-1,0,0,1,0,0,1,-2,-1,0,-1,0,0,2,-1,-2,-1,1,0,0,-2,1,0,1,0,-1,1,-1,1,-1,-1,-1,1,1,1,-1,1};
			381: counter1_out = '{0,1,1,-1,1,0,0,-2,-2,0,1,-3,0,0,1,-1,1,1,-1,0,0,1,0,0,-1,-1,-4,1,1,-2,-1,1,-2,-1,-1,0,2,-3,0,1,1,1,1,1,-1,-1,0,-1,1,0,1,-3,-2,0,0,1,-1,0,1,-1,-1,-1,1,-3,0,-2,0,-1,1,0,0,-1,0,-1,-2,0,0,0,0,-1,0,0,-1,1,1,2,1,0,-1,-1,0,0,-2,0,2,0,0,1,0,-1};
			382: counter1_out = '{1,0,1,0,1,0,-1,-1,-1,1,-1,0,-2,2,0,0,0,0,-1,1,0,1,0,0,1,1,0,3,1,0,1,-1,-1,0,0,0,1,-2,1,0,-1,-1,-1,-1,-1,-2,0,-1,0,1,2,0,0,1,0,0,0,0,0,0,1,1,0,-1,1,-1,0,0,-1,2,0,-2,-2,0,0,-2,1,1,0,0,-1,1,1,-3,1,0,0,1,0,0,-2,0,-2,0,-2,0,0,0,-1,-1};
			383: counter1_out = '{1,2,0,0,0,-1,-1,-1,-2,1,-1,0,0,0,2,1,1,0,-1,2,0,0,0,0,0,0,2,1,-1,1,0,0,-1,-1,-1,-2,2,-2,1,-1,-1,0,-1,0,-3,0,1,-2,0,-1,-2,2,0,-1,0,-1,-1,1,0,-2,2,-1,1,1,-1,1,1,-1,1,-1,0,0,-1,-1,-1,2,0,-2,0,-1,-1,0,0,-1,0,1,-1,1,1,-2,-1,0,0,0,-2,1,1,1,1,-1};
			384: counter1_out = '{0,-2,0,1,0,1,-1,0,-1,0,2,0,-2,0,0,1,-2,0,-1,1,0,1,0,0,0,1,1,-1,2,2,0,0,-2,-1,1,-1,0,-1,0,-1,0,0,0,-1,1,-1,1,-1,-2,-1,0,1,1,1,-1,-2,-2,-1,2,-1,-2,1,0,-1,-1,0,1,0,3,0,-1,-1,2,-1,0,0,1,-2,1,-1,-2,1,-1,-1,1,1,-2,-1,0,-2,-2,1,1,-3,1,0,-1,1,-2,1};
			385: counter1_out = '{0,-2,2,-1,-2,0,-2,-1,-1,-1,0,0,1,1,-2,-1,0,-1,1,2,-1,2,1,2,-1,1,1,-2,-1,0,-1,0,-1,0,1,-2,1,0,0,-2,-1,1,1,-1,1,-1,-1,0,0,1,0,-1,-2,-2,-1,-1,-1,2,1,0,0,1,1,1,0,1,1,0,2,0,1,1,1,-1,-1,2,-2,0,-1,-1,-1,1,-2,-1,3,2,-2,-1,1,-2,-3,0,-1,1,-1,1,0,1,0,-1};
			386: counter1_out = '{-1,2,1,-1,-1,1,1,0,0,0,0,1,2,0,0,-2,1,0,0,2,2,0,1,0,-3,0,0,-1,1,-1,0,1,-1,-2,1,-1,1,-2,0,-3,0,1,0,0,0,-3,-1,0,0,-2,-1,1,-1,0,-1,-1,0,0,0,2,1,1,-1,0,0,1,-1,1,1,0,-1,-1,-2,2,2,2,-1,0,1,0,-3,1,0,0,1,2,-1,-1,-2,-1,-1,0,1,1,-3,1,0,0,-1,0};
			387: counter1_out = '{0,-3,-1,1,-1,-1,0,-1,-2,-1,0,-1,0,2,-1,-1,0,1,-1,1,-2,-2,1,0,0,2,0,-1,-1,0,1,0,0,0,1,0,1,-2,1,1,-1,-1,0,0,1,-1,3,1,0,-1,-1,1,0,-1,-1,0,-1,-1,-1,-1,0,1,0,0,0,0,0,0,1,2,-1,0,1,2,1,1,-2,0,0,1,0,1,0,0,1,-1,-1,1,0,-1,0,0,-1,1,-1,3,1,1,1,1};
			388: counter1_out = '{1,1,0,0,1,2,-1,0,-1,1,0,0,0,-1,1,1,2,-1,0,0,1,0,1,-1,0,2,0,-1,-2,1,0,-1,0,1,2,1,-1,0,1,-1,-1,-1,-1,0,0,0,-1,-1,0,3,1,0,1,0,-1,0,0,0,-1,0,0,0,3,-1,2,-1,-1,2,1,-1,0,1,-2,0,1,1,-2,-1,-1,0,-1,-2,-1,0,1,0,1,0,1,-2,1,0,-2,0,1,0,0,0,-3,1};
			389: counter1_out = '{1,0,0,-1,0,-1,2,-1,0,0,0,-1,1,-1,-1,-1,-1,-1,-1,0,-1,1,1,-1,0,0,0,1,1,1,0,2,1,-1,0,0,1,-1,1,1,0,-1,-1,0,0,1,1,-3,-1,-1,-1,-1,2,-2,0,1,1,1,-1,-2,1,-1,0,0,-2,-1,-2,-1,0,0,1,-2,1,-2,0,0,-1,1,-1,2,-1,0,0,0,2,-1,-2,0,0,-1,2,-1,0,1,0,-1,1,-1,-1,1};
			390: counter1_out = '{-1,0,0,1,-1,0,2,1,1,0,-1,1,0,0,0,1,1,1,-1,-1,0,1,-1,-1,0,1,1,-1,0,0,-1,0,0,-2,1,1,0,1,1,-1,2,1,-1,-1,0,0,-1,1,-1,0,-1,-1,0,1,0,1,0,-1,0,1,1,2,0,-1,-3,1,0,0,0,0,0,1,-1,1,-1,1,2,-1,0,1,0,1,1,0,0,1,-1,0,1,-1,-2,0,-2,0,-1,0,0,0,0,1};
			391: counter1_out = '{1,1,1,1,0,0,0,-1,0,0,-1,0,-1,-1,0,0,2,0,0,0,1,-1,0,1,-1,-2,1,1,-1,0,0,1,-1,1,1,2,-2,-1,0,0,1,-2,1,0,0,0,0,-1,-2,-1,-1,0,2,-3,1,-1,0,0,1,0,0,0,1,1,0,-1,0,-2,1,2,0,-1,-2,0,1,-2,1,1,0,-1,-1,1,0,0,-1,1,0,0,0,0,2,0,-2,1,-1,-1,0,-1,0,-2};
			392: counter1_out = '{-1,1,2,0,0,0,0,0,0,0,-1,1,0,0,1,0,0,0,1,-1,0,0,1,0,0,0,1,-1,0,1,-1,-1,0,-1,0,1,0,0,-2,-2,0,0,2,-1,0,0,-1,-1,0,0,-1,-1,0,1,1,0,0,0,0,0,-1,0,0,0,0,0,0,3,2,1,0,-1,0,1,1,0,-1,1,1,0,1,0,0,-1,-1,0,1,1,0,-1,1,0,-2,-1,0,0,0,-1,0,1};
			393: counter1_out = '{2,0,0,0,-2,-1,-2,0,0,0,0,0,2,0,0,0,0,0,0,0,0,0,0,0,0,-2,-1,2,0,-1,2,0,-2,-1,0,1,0,0,-2,2,1,0,-1,1,1,1,0,-1,-1,0,-1,0,-1,1,0,0,1,-1,0,0,-1,0,0,0,1,-1,-1,0,0,3,1,1,0,1,0,1,-1,1,1,-1,0,2,0,1,1,0,1,1,0,-1,0,2,1,1,1,1,1,0,0,1};
			394: counter1_out = '{0,-2,-1,1,0,0,0,0,-1,0,1,0,3,-1,-1,2,1,2,-1,1,-1,0,1,-2,0,2,1,1,-1,0,-1,-1,1,1,-3,0,0,0,2,-1,1,0,0,0,-1,-1,0,0,-1,0,-1,0,0,0,0,2,0,-1,-1,0,0,-1,2,1,0,-1,0,0,-1,1,0,0,0,0,0,-1,-1,2,-1,0,1,-1,1,-1,-1,0,1,-1,0,1,-1,0,0,1,-1,1,-1,2,2,1};
			395: counter1_out = '{0,0,-2,1,1,1,0,-1,-1,-1,0,-1,0,-2,-1,-1,-1,2,0,1,-1,2,1,-2,-2,1,0,1,0,-2,-1,0,0,0,0,1,-1,1,0,1,-1,0,-2,-1,-1,1,3,2,0,-1,0,-1,1,1,1,1,0,1,1,1,3,1,0,1,-2,0,1,0,1,0,-1,-2,-1,-1,0,-1,-1,1,-1,-1,-1,0,0,1,1,1,0,2,0,1,1,0,3,-1,1,1,1,2,-1,1};
			396: counter1_out = '{-2,0,2,-2,1,-1,2,-1,0,3,0,1,2,-1,0,-2,1,0,-1,1,-2,0,0,-2,0,-1,-1,0,-1,-3,-1,1,0,-1,0,0,1,0,0,0,0,0,-1,0,0,1,0,0,-1,0,0,2,1,1,0,0,1,1,1,1,2,2,-1,1,-1,2,0,0,2,0,0,1,-1,2,-1,0,0,-1,0,-2,0,2,-1,0,-2,-1,-1,-1,0,0,0,0,0,0,0,0,-1,0,-1,-1};
			397: counter1_out = '{0,0,0,-1,1,-1,-1,-1,-1,-2,-2,0,-1,0,-2,-1,1,1,-1,1,-1,2,0,0,2,0,0,1,2,0,1,0,-2,0,0,0,-1,1,1,-1,0,1,2,0,0,0,0,0,1,-3,0,1,0,-1,2,1,0,-2,0,1,0,3,0,0,-1,-2,0,-1,2,0,-1,2,-1,0,1,-2,-1,1,-2,1,-1,0,1,0,1,0,-2,-1,-1,1,0,1,1,-1,3,1,-2,1,0,0};
			398: counter1_out = '{1,-1,1,-1,-1,1,0,-2,0,-1,1,1,0,0,0,1,0,1,0,-1,-1,0,0,0,-1,-1,1,1,1,1,-1,1,0,0,-1,-1,0,0,-1,0,2,1,0,0,1,1,-1,-1,-1,-3,-1,-1,-1,0,-1,0,-2,0,0,-1,2,1,-1,1,0,-1,0,0,1,0,0,-1,1,1,1,2,-3,0,-1,2,0,2,0,-2,1,0,-2,1,-1,0,0,0,1,1,0,0,0,1,-1,-1};
			399: counter1_out = '{-1,0,2,-1,1,-2,0,0,0,1,-1,0,0,-1,-1,-1,1,1,0,-1,-1,1,0,2,0,0,0,0,0,-1,-1,-1,-1,1,-4,-1,1,0,-2,-1,1,2,0,0,1,-2,0,0,1,-2,-1,1,-1,-1,1,1,0,0,0,1,0,0,-1,2,2,3,-1,0,2,0,0,0,0,0,1,-1,0,-1,-2,0,1,2,-1,-1,0,1,0,3,-1,-1,1,1,2,2,0,2,1,0,0,0};
			400: counter1_out = '{0,1,1,-1,0,-3,1,0,0,2,-1,-1,-1,-2,1,0,0,1,-1,0,0,0,0,0,2,0,0,1,0,1,0,-1,-1,1,0,0,0,1,0,-2,0,2,1,-1,1,-1,-1,-1,0,-2,0,0,0,-1,0,-1,-1,2,0,0,0,2,0,0,1,-1,1,0,-1,0,1,1,1,0,0,2,0,2,-1,0,1,2,1,0,2,2,-2,-1,-1,-1,0,0,0,1,2,-1,1,0,-1,-1};
			401: counter1_out = '{0,1,0,0,0,0,-1,1,2,0,-2,0,0,0,0,-1,-2,2,1,0,0,0,0,-1,-2,0,0,0,1,-1,0,-1,3,1,1,0,-1,-1,1,-1,-1,1,1,1,0,-1,-2,0,0,-1,1,2,0,1,0,1,-2,0,1,0,-1,1,0,0,-1,0,0,1,-1,0,-2,1,0,1,0,1,0,1,1,1,-1,0,-1,-1,0,0,-1,0,-1,1,-1,-1,-1,3,1,-2,0,0,1,0};
			402: counter1_out = '{-1,0,0,-1,-3,0,0,1,-1,0,0,-2,-1,0,0,0,-1,1,0,-3,0,0,-1,0,-2,-1,2,1,1,2,1,0,-2,1,-1,-1,-1,-2,0,-1,0,-1,2,-1,-1,0,-2,0,0,-1,-2,1,1,0,1,1,0,1,-1,1,0,2,-1,0,0,-2,1,0,1,-1,2,1,0,0,-1,0,-2,1,1,0,1,2,-1,-1,0,0,0,-1,-1,0,0,1,1,2,1,0,-2,0,0,0};
			403: counter1_out = '{1,-1,0,2,-1,0,-1,-3,0,0,1,-2,0,2,1,0,-2,-1,1,0,-1,-1,1,4,0,1,0,-1,1,0,1,1,-1,1,-1,-1,0,0,3,-1,1,2,1,1,0,-3,-1,0,-1,-1,0,0,0,0,2,0,1,0,1,0,0,3,0,1,0,-2,0,1,-2,-1,0,2,-2,-1,2,0,2,0,2,-1,0,2,-2,0,-2,1,-1,1,0,2,0,0,1,-1,-2,0,-1,3,-1,0};
			404: counter1_out = '{2,0,1,2,1,0,1,-2,-1,0,0,-2,-1,0,1,1,-1,-1,-2,0,-1,-1,1,0,0,0,1,-1,2,1,2,-1,0,0,1,-1,-1,-1,0,2,0,2,0,-1,-1,-1,-2,1,0,-1,-1,1,2,0,1,3,0,-1,1,0,-1,-1,-1,1,1,-1,1,-1,0,0,0,1,-1,-4,1,1,0,1,1,0,0,1,-2,0,0,0,0,0,2,0,1,1,2,3,-2,0,-2,0,-3,0};
			405: counter1_out = '{4,0,2,0,-1,-1,1,0,0,1,2,-1,0,-2,0,-1,0,-2,0,0,0,-1,1,0,0,2,-1,1,-1,1,1,2,-2,0,0,1,2,1,0,0,-1,0,-1,0,-1,-1,-2,-2,0,-1,0,-2,-2,1,-1,1,0,-2,0,-1,-1,-2,1,0,0,1,-1,-1,0,1,-1,0,1,-1,0,2,1,-1,-1,0,0,-1,-2,-1,0,-1,-1,-1,-1,0,0,0,0,-1,-3,0,-1,0,-2,-1};
			406: counter1_out = '{2,0,0,1,0,0,1,0,1,1,-1,-1,0,1,2,-1,0,-1,0,-1,0,0,0,0,1,0,0,1,1,-3,0,0,1,0,2,0,0,-1,2,-1,-1,-1,-1,0,0,2,-2,0,2,0,1,-2,1,1,1,1,-1,-2,-2,1,-1,-1,-1,1,0,-1,1,0,0,2,2,1,-1,1,1,0,3,1,0,-1,0,0,-2,1,-3,1,0,-1,1,2,-1,0,-1,0,-1,1,1,-1,-2,-1};
			407: counter1_out = '{1,1,0,1,0,0,-1,0,2,-1,-1,-2,-2,-1,-1,-1,2,1,-1,0,0,1,0,-1,3,0,-1,1,0,-2,-1,1,0,0,0,1,1,2,-1,-1,1,-3,0,1,0,-1,0,-1,1,0,0,-2,-2,1,-1,1,1,0,1,-1,0,0,1,0,2,0,1,-1,1,-1,3,-1,-1,-2,0,1,2,-1,0,-1,-2,0,-3,1,1,0,0,1,2,-1,0,2,0,0,1,0,1,-1,1,0};
			408: counter1_out = '{-1,-2,2,-1,2,-1,0,-1,-1,-1,0,-2,-1,1,3,1,0,-1,1,-1,0,0,-2,0,-1,0,-2,2,0,-1,0,1,0,-1,-1,1,1,0,-1,1,0,-2,0,0,-1,1,1,-1,0,-1,0,-3,0,1,1,0,1,1,0,-2,-1,0,-1,-1,1,0,0,1,0,0,1,0,1,0,-1,2,2,0,0,-1,1,-1,-3,-1,2,1,0,-1,0,1,-1,0,-2,-1,-3,1,2,2,-1,0};
			409: counter1_out = '{0,-2,2,0,1,-1,-1,-1,1,0,-1,-2,0,0,1,-1,1,-1,0,0,0,1,0,0,2,1,1,1,-1,-1,-2,-2,0,1,0,-1,-1,-2,1,-1,-2,0,-2,0,0,1,0,0,-1,-1,0,-2,1,2,1,1,0,0,1,-1,1,1,1,-1,1,-1,2,-1,1,0,-1,0,0,0,-1,-1,-1,0,-1,0,0,-1,-1,-1,-1,2,0,0,0,0,-2,1,1,-1,0,-1,0,-1,-2,-2};
			410: counter1_out = '{0,0,4,-2,1,0,1,1,-1,-1,0,0,0,1,-1,0,1,-1,-1,2,-1,2,0,0,0,-1,0,0,0,-1,0,1,0,0,1,-2,1,-1,-1,1,0,-1,1,-2,1,0,-1,0,0,0,-1,0,0,0,-1,-1,-1,1,1,0,0,1,0,0,1,-1,3,-1,1,0,1,1,-1,0,0,0,-1,-1,-2,-1,1,-1,-1,0,-1,1,1,0,-1,0,-1,0,0,0,0,1,0,0,-1,1};
			411: counter1_out = '{0,0,2,2,0,-1,-1,0,-1,1,1,-2,-1,1,1,1,-1,0,-1,1,0,0,0,2,-1,0,0,0,0,0,1,0,1,0,-1,-1,2,-2,-1,-1,0,-1,-1,-1,1,-1,-3,0,1,1,-1,-2,3,2,0,0,1,1,-1,1,2,1,-1,0,1,0,0,0,0,-2,-1,0,-1,-1,0,1,0,1,-1,-2,-2,1,1,-1,-1,2,1,1,1,0,-1,0,-1,0,0,0,-1,-1,0,-2};
			412: counter1_out = '{-1,0,1,0,1,1,1,-1,1,-1,-2,-2,1,1,-1,0,-1,0,0,0,0,0,0,0,1,0,1,0,0,-2,-1,0,-1,1,1,-1,0,-2,1,1,-1,2,-1,1,0,0,-1,0,0,0,1,1,0,0,0,-1,0,2,0,1,2,0,0,-1,0,1,0,0,3,-1,0,0,0,0,-3,0,-1,-1,0,1,0,1,-1,1,1,1,2,0,-3,0,-2,-1,0,2,0,1,-1,-1,-1,0};
			413: counter1_out = '{-1,0,2,0,-1,0,0,-1,1,-1,-2,0,1,-1,1,-1,-1,1,3,0,1,0,0,1,0,0,0,0,0,-1,0,-1,1,0,-1,0,2,-3,-1,-1,-1,0,0,0,-1,1,0,-1,1,0,1,0,-1,-1,-3,2,0,-1,0,1,1,0,1,-1,-1,1,0,-1,1,0,0,-2,-1,3,-1,0,0,0,1,-1,0,-1,0,1,1,-1,0,0,-1,-1,-1,0,-1,0,0,1,0,1,0,0};
			414: counter1_out = '{1,0,2,0,-2,-1,-2,0,0,0,1,-1,-1,0,1,1,0,1,0,0,0,0,-1,0,-1,0,1,-1,1,2,-2,-1,-1,0,1,1,0,-1,-1,1,0,-1,2,0,1,0,-1,0,-1,1,-1,3,-1,0,0,0,-3,0,1,-1,1,0,0,0,1,-1,-2,0,0,0,0,1,1,2,1,0,0,0,-2,0,1,1,-1,-1,1,0,1,0,0,-2,-1,1,0,2,-1,1,-1,0,-1,0};
			415: counter1_out = '{-2,0,0,-1,0,0,0,3,-1,1,0,0,-1,-1,0,-1,-1,-1,-1,-1,-1,-2,-1,0,0,0,-1,1,1,0,-1,-1,0,0,1,1,0,-1,0,-1,-1,-2,1,0,0,0,1,1,2,-1,-2,0,-1,0,-1,0,1,0,1,-3,-1,0,0,1,1,1,1,-1,2,-1,2,-1,-1,1,2,0,0,0,-1,0,0,-2,0,0,0,-1,-2,-1,0,0,-1,0,0,1,0,0,0,-1,0,1};
			416: counter1_out = '{2,-1,1,0,1,-1,1,1,-2,1,0,1,1,0,-1,0,0,1,2,1,1,-1,0,0,0,0,2,2,-1,2,1,-1,1,-1,0,0,-1,-1,-1,0,1,0,1,-1,0,1,0,0,1,0,1,1,-1,1,0,-1,1,2,0,1,2,2,0,-1,1,1,-1,2,1,0,2,0,-1,1,2,-1,-2,-1,-2,1,1,0,0,1,0,-1,1,-2,2,0,-2,1,-1,1,1,0,-1,-1,-1,0};
			417: counter1_out = '{1,-1,0,0,1,2,1,0,3,0,0,-1,0,0,-1,1,-1,2,-1,-1,0,0,1,0,0,-1,0,-1,0,-1,-1,2,1,1,1,0,0,0,1,0,-1,-1,1,-1,-1,0,-1,1,-1,0,0,-1,1,0,-2,2,0,1,1,2,0,0,0,0,0,0,0,1,-1,0,-1,1,0,-1,-1,-1,-1,0,0,1,0,0,1,1,1,-1,-1,0,1,-1,-1,-1,0,0,-1,1,-1,0,1,0};
			418: counter1_out = '{1,0,1,1,1,0,2,-1,0,0,0,1,-1,1,-2,0,0,0,-1,0,1,1,0,0,2,1,-1,0,-1,0,-1,-1,0,0,1,-1,1,1,1,-1,-2,0,1,-1,-1,0,0,1,1,0,1,2,1,0,-1,-1,0,1,1,3,1,0,1,0,0,0,0,1,-1,1,2,-1,0,0,2,-1,0,0,-2,0,0,-1,1,1,1,1,0,1,-1,-1,-1,-1,1,1,0,-2,0,2,0,1};
			419: counter1_out = '{0,-2,-1,2,-2,0,-1,1,1,1,0,0,-1,1,-1,0,1,3,2,1,0,0,1,-1,-1,2,-1,-1,-1,0,1,0,1,0,0,-1,0,2,-1,1,-1,-1,1,0,0,1,0,-2,-2,1,0,0,0,0,0,0,0,0,1,1,0,1,1,1,-2,1,1,-2,1,1,1,0,0,2,1,0,-1,1,-1,-1,0,0,0,0,-1,1,0,-1,-1,-1,-1,1,2,1,0,0,0,-1,1,0};
			420: counter1_out = '{1,0,0,0,0,1,0,-1,1,0,1,1,0,0,2,1,1,0,1,-1,-2,1,-1,0,1,-1,0,1,-2,-2,2,1,-1,0,0,0,0,1,1,-2,-1,3,1,0,0,0,-1,-1,1,0,1,-2,-1,-1,0,1,0,0,-1,0,-1,0,-1,-1,-1,2,0,0,0,1,0,-1,0,-1,2,1,-1,0,-1,-2,1,1,0,1,1,0,0,0,-1,0,1,2,0,0,-2,1,0,-1,0,0};
			421: counter1_out = '{0,1,0,-1,0,0,0,-1,-1,0,0,0,-2,-1,0,1,0,-1,-1,0,0,1,0,-2,-1,-1,0,2,2,1,-1,1,-1,-2,2,-1,1,0,1,-1,-2,0,0,-1,-1,0,0,-2,0,0,0,0,0,-1,0,1,0,0,0,0,1,1,1,1,-1,2,0,0,3,1,-1,1,1,1,0,1,2,0,0,0,0,-1,1,0,0,-1,-1,-2,0,1,-1,-1,0,0,0,0,0,-1,1,0};
			422: counter1_out = '{0,2,0,-2,0,-1,0,-1,1,0,1,0,0,1,0,0,1,1,-1,-1,1,0,-1,1,0,-2,2,1,0,-1,0,0,0,1,1,0,-3,0,-1,-2,1,0,1,-1,-1,1,-1,-1,-1,1,1,0,1,1,0,0,0,-1,0,1,1,0,0,0,0,-1,0,0,-2,1,2,-2,1,0,2,2,1,1,0,0,0,-1,1,0,1,0,0,0,1,0,0,-1,0,2,-1,1,0,-1,2,-2};
			423: counter1_out = '{-1,2,0,-2,2,-1,0,-2,1,0,0,0,-1,-1,1,1,0,0,0,-2,0,0,0,1,0,0,-2,0,-1,-2,0,-1,-2,-1,0,0,0,-1,-1,1,-2,-1,-1,-1,-1,0,0,2,-1,0,0,0,0,0,-1,-1,0,1,1,-1,-1,2,-1,1,0,0,1,-2,-1,0,0,-2,0,-1,0,-1,0,0,0,1,-1,2,0,1,0,2,-1,-1,1,1,-1,1,0,1,0,1,-1,0,0,0};
			424: counter1_out = '{0,0,0,0,1,2,1,0,0,-1,0,0,1,0,-1,1,0,-1,-1,-1,-1,0,1,-2,-2,1,0,0,0,1,0,2,1,-1,0,0,2,1,0,1,1,0,0,-2,0,0,-1,0,0,1,-1,1,-2,0,0,2,1,0,0,1,-1,0,0,1,1,1,0,1,0,1,0,-1,-1,0,0,0,-2,0,-1,-1,-1,0,-1,-2,1,1,-1,0,-2,1,0,0,-1,2,-1,0,-2,-1,0,1};
			425: counter1_out = '{0,1,1,0,0,-1,-1,-1,0,-1,1,3,0,-2,-1,-1,0,1,0,0,0,0,0,1,-1,1,1,0,1,0,-1,0,3,-1,0,2,0,-1,0,0,-1,-2,-1,2,0,-2,0,-3,-1,-2,-2,0,-1,0,1,1,-1,0,0,1,1,2,0,1,-1,2,0,1,-1,-1,0,-1,0,1,1,-1,-2,-1,0,3,1,-1,-1,-1,-1,0,-2,-1,-2,1,-1,0,0,1,0,0,2,-1,0,2};
			426: counter1_out = '{1,0,0,-1,-1,0,0,2,0,-2,0,0,1,0,1,0,-2,2,-1,1,-1,1,1,0,-1,0,3,0,0,1,-2,0,1,0,-2,-1,-2,-2,0,0,0,-1,0,1,0,-1,0,2,-2,-5,0,0,1,-2,-1,0,0,1,1,0,0,0,1,0,0,0,1,1,0,-1,-2,2,0,0,0,1,-3,-1,0,0,-1,-1,0,1,1,2,-1,0,0,-2,3,1,1,0,0,1,0,0,2,1};
			427: counter1_out = '{1,0,1,-2,-2,0,-1,0,1,1,0,-1,0,0,1,0,0,1,-1,0,2,0,1,0,0,-1,0,2,1,-1,-1,0,0,1,-2,0,0,-1,2,-1,1,1,1,0,0,0,-1,-1,-1,-5,0,0,-1,1,0,1,-1,0,1,-1,0,2,-1,2,3,0,0,1,0,-2,0,1,0,2,-1,2,-2,0,-2,2,1,1,0,1,-1,-2,0,0,0,0,2,-1,0,2,1,1,1,1,0,1};
			428: counter1_out = '{1,1,2,0,-1,0,0,0,-3,1,-1,-1,1,0,1,0,0,0,-1,-1,-1,0,1,0,-1,1,1,0,2,0,-1,-2,-1,1,0,0,-1,0,-1,1,-1,1,1,2,2,0,-2,0,-1,-5,-2,0,1,0,1,0,-1,0,0,0,0,1,-2,-1,-1,-1,0,0,1,-3,1,0,0,1,0,0,-1,2,1,1,0,0,0,-1,0,0,0,-1,-1,1,0,0,1,2,-1,0,-1,1,2,0};
			429: counter1_out = '{2,-2,0,1,0,-2,1,-1,-1,0,0,-1,-1,0,-1,1,-1,0,0,0,1,1,0,1,0,0,1,0,1,-1,-1,0,1,-2,0,0,-2,-1,-2,-1,-1,0,-1,2,1,-1,-1,0,0,-2,-1,0,0,-1,0,1,-2,1,-1,-1,-2,1,0,0,0,-1,1,0,-2,-1,1,1,1,-1,-2,1,-1,0,1,-1,0,0,0,0,0,-1,-1,2,-1,-2,0,-1,-1,2,-1,-1,1,0,0,1};
			430: counter1_out = '{1,-1,1,-1,-1,1,1,-3,-1,-1,1,-1,0,0,1,0,-1,-1,0,-2,1,2,0,1,-1,0,1,0,0,0,0,0,0,1,-1,-3,1,1,0,-2,-1,0,0,1,1,-1,-1,-2,2,-2,-2,0,0,0,1,-1,-1,0,1,1,1,3,1,2,1,0,-1,-1,1,1,0,0,-2,-1,-1,0,-1,-1,0,0,-1,0,-1,1,2,-1,0,-2,2,1,-1,-1,-1,1,0,0,0,0,-1,0};
			431: counter1_out = '{2,-1,0,-2,-1,1,0,-3,1,-1,1,0,1,1,0,1,0,1,0,0,0,1,-1,-1,0,-1,0,2,0,0,0,0,2,0,1,-1,2,-2,0,-3,-1,2,-2,1,0,-1,-1,0,-2,-1,-2,-1,1,-2,-2,0,-2,1,-1,0,2,0,0,-2,0,0,-1,-1,-2,0,1,0,-1,-2,0,-1,1,-1,0,0,0,-1,-1,0,1,0,0,0,1,1,1,-1,-1,2,-1,1,1,0,-1,1};
			432: counter1_out = '{2,-1,-2,0,-2,-1,1,0,1,1,1,-1,0,-1,3,0,0,0,1,0,-1,0,-1,-1,2,-2,0,-1,2,0,1,2,-2,-1,0,2,0,0,2,-2,0,2,1,0,1,0,-1,1,1,0,0,0,1,-1,-1,2,0,0,2,0,0,-3,2,-1,0,-2,1,0,1,0,1,0,1,-2,0,1,-1,1,0,-1,1,1,0,2,1,0,-1,0,0,0,2,0,0,1,-2,-1,-2,2,0,1};
			433: counter1_out = '{2,0,-1,0,2,-2,0,-1,-1,0,1,-1,0,-2,0,0,0,-1,1,1,-1,1,0,-1,0,0,-1,0,0,0,-1,-1,1,1,2,1,0,1,-1,-1,-3,1,0,0,0,0,-2,0,-1,-1,-1,-1,-2,-1,-1,2,0,1,0,-1,-2,-1,1,0,-1,-1,-2,-2,0,0,2,0,0,1,1,0,2,1,-1,-1,0,2,0,-2,1,-1,-1,1,0,3,1,0,-2,-1,-3,-1,-1,1,-2,0};
			434: counter1_out = '{0,-1,3,0,0,0,0,1,0,2,-1,-2,-1,1,0,0,0,-1,1,2,0,-1,0,0,2,2,-1,0,0,-1,3,2,0,-1,3,1,-1,-1,0,-1,-3,1,-2,0,-2,-2,1,0,1,0,1,-2,0,-1,0,1,0,0,-4,-1,0,1,1,2,1,0,0,0,1,0,0,0,1,1,0,1,1,0,-2,-4,-1,1,-1,0,0,1,0,1,1,1,0,2,0,-1,-2,0,0,1,0,0};
			435: counter1_out = '{1,-1,0,1,0,-1,1,-1,2,0,1,-1,-3,-2,-1,0,-1,1,0,-1,1,2,0,-1,1,1,-3,1,0,0,2,0,2,0,0,1,1,1,1,-1,0,-1,-1,2,1,-1,1,1,-1,-1,-1,-2,1,0,0,1,1,2,0,-1,0,-1,-2,0,1,-2,0,-2,0,-1,0,2,-1,0,-2,0,1,0,-1,0,0,3,-1,-1,1,-1,-1,-1,1,-1,-2,1,-2,1,-1,-3,0,0,-1,0};
			436: counter1_out = '{2,1,2,1,0,-1,0,-1,0,-1,0,-2,-3,2,0,0,0,-2,0,-1,0,0,0,-2,1,-1,0,0,-1,-1,-2,-1,0,2,0,0,2,0,-1,0,-1,1,0,0,3,0,-1,-2,1,-1,0,-2,0,1,0,0,-1,0,2,0,1,1,-1,1,1,-1,0,-1,1,-1,0,-1,0,1,0,1,1,1,-3,-2,0,1,-1,-1,0,-1,1,0,0,0,-2,1,0,0,0,0,-1,0,0,-2};
			437: counter1_out = '{0,1,1,-2,0,-2,1,-1,-1,2,0,-2,0,1,-1,1,0,0,-3,1,-1,1,0,2,1,-1,-2,0,1,1,0,1,0,-1,-1,-1,1,0,0,0,1,-1,-1,-1,-2,1,2,-2,0,0,1,-2,1,1,0,1,0,1,3,-2,1,1,0,1,0,-3,1,1,1,-1,0,0,0,0,1,0,-1,1,-2,1,-1,1,-1,0,0,1,-1,1,0,0,0,0,0,0,0,-1,1,-1,-1,0};
			438: counter1_out = '{1,0,0,-1,1,1,0,-2,0,0,1,-1,-1,2,0,0,-1,-2,-1,1,0,1,1,2,1,1,2,0,1,0,0,-1,0,0,0,-2,2,0,1,0,0,1,0,-1,2,0,1,0,1,1,0,0,1,0,-1,2,0,2,0,-1,3,-1,-1,2,0,0,0,0,1,0,2,-1,0,1,-2,2,-2,2,1,1,0,1,-2,-1,0,1,0,1,-1,0,-1,0,1,0,1,-3,-1,-1,3,1};
			439: counter1_out = '{1,1,3,1,0,-1,1,-2,0,0,0,0,1,0,0,0,-1,0,1,1,-1,2,-1,0,-1,-1,1,0,-1,0,0,-1,0,0,2,-4,1,-2,1,2,-1,-1,0,-1,-1,0,0,0,-1,-2,1,0,0,0,0,-1,-1,0,0,2,0,1,0,0,0,1,-1,0,1,0,1,-1,1,2,2,1,0,0,2,2,0,-1,1,1,1,-2,-1,1,1,1,-1,1,-1,-1,0,0,-1,-1,-1,0};
			440: counter1_out = '{1,2,1,-1,0,0,0,1,0,-2,-2,1,0,-1,0,-2,-1,0,-1,0,-2,0,2,0,-1,1,0,-1,1,0,-1,-1,0,0,-2,0,0,-1,-1,-2,-1,0,1,-1,-1,1,1,-2,2,-1,1,0,-1,1,-1,0,0,0,-1,1,1,1,0,0,1,1,0,1,-1,1,0,1,1,2,0,0,-1,2,-1,0,0,-1,0,-1,1,0,0,1,-2,0,-1,1,-1,0,0,0,-1,0,2,1};
			441: counter1_out = '{0,-2,2,0,0,2,-1,1,0,1,-1,1,-2,1,0,0,0,-1,1,0,1,0,0,-1,0,0,-2,-1,0,-1,-2,-2,1,1,1,0,-1,0,1,-1,2,-1,0,-1,-1,-3,1,0,2,1,0,-2,0,-1,0,0,-2,0,-1,1,1,0,0,3,2,2,-1,0,1,0,-1,0,-1,2,2,1,0,0,0,0,-1,-1,1,1,-2,2,-1,-1,1,0,0,0,1,1,-1,2,-2,-1,0,-1};
			442: counter1_out = '{0,0,2,1,-1,1,-1,-1,0,0,0,-1,-1,1,1,-1,1,-1,0,2,0,1,0,1,0,1,-2,-2,-2,0,0,-1,0,0,1,0,-1,-4,2,-1,1,1,0,-1,-1,-1,0,-1,1,-2,0,0,-1,0,-1,1,-2,2,1,0,0,1,0,-1,0,2,0,2,1,1,3,0,0,1,2,1,-1,2,1,0,0,0,-1,1,0,1,-2,0,-1,-1,0,0,-2,1,-1,0,0,-1,1,0};
			443: counter1_out = '{1,-1,0,0,0,1,0,-1,-1,1,-2,0,0,-1,2,1,0,0,-1,-1,-1,1,0,0,-1,0,-1,0,0,1,2,-1,-1,-1,3,-1,1,0,0,-2,0,0,1,-2,-2,-1,0,2,1,0,-2,0,0,1,0,0,-2,1,1,-1,1,4,0,1,0,0,1,-1,1,2,2,1,0,2,1,1,-1,0,3,1,0,1,2,0,2,-3,-1,1,1,0,-1,-2,0,0,-1,-1,-1,0,1,0};
			444: counter1_out = '{-2,1,-1,-2,-1,0,-1,2,0,1,-1,2,2,0,1,0,0,0,1,0,0,1,-2,0,0,0,-1,1,0,2,3,-1,-1,1,-1,2,1,0,-1,-1,-1,-1,0,-1,1,0,0,-1,1,0,2,0,1,0,0,-1,-1,0,0,-1,2,0,0,0,1,0,-2,1,-2,2,-1,-1,-1,-1,2,2,1,0,-2,-1,0,-2,1,0,0,-1,0,-2,-1,0,1,0,1,0,0,-1,2,0,-1,-1};
			445: counter1_out = '{-1,0,-2,0,0,1,-1,0,0,1,-1,-1,0,0,-1,0,0,0,0,2,-1,0,-1,1,0,-2,-1,0,1,1,2,1,-1,0,1,0,2,2,0,3,-1,0,-1,1,1,0,1,0,-3,-1,-2,1,1,2,0,-1,0,1,-2,0,0,-1,-1,1,-1,0,-1,-1,0,0,-2,0,1,1,0,-1,-1,1,-1,-1,1,1,0,0,0,0,0,-1,0,0,-1,0,0,1,0,0,1,0,-1,2};
			446: counter1_out = '{2,-1,-2,2,0,-1,1,0,0,1,0,2,-1,0,0,0,-1,-1,-2,0,0,0,1,0,1,0,-2,1,1,1,0,1,2,-1,1,-1,0,-1,2,1,-1,-1,-1,0,0,-1,-1,0,0,-1,-1,1,0,2,-1,-1,0,-1,0,0,0,2,1,-1,1,1,0,-1,1,-1,-1,0,0,-1,0,1,-2,0,0,-1,-1,-1,0,1,1,-2,-2,0,1,-1,-2,0,1,0,-1,0,2,0,0,-1};
			447: counter1_out = '{0,-1,-3,1,2,2,2,-1,0,0,-1,2,0,0,-1,0,2,0,-1,1,-2,0,1,-1,0,0,-1,-1,1,-2,-2,0,-1,1,-1,2,0,-2,1,1,2,-2,-2,0,2,-2,1,0,1,-1,-1,0,0,0,0,-1,0,0,-1,0,-1,0,0,-1,1,0,1,0,1,1,0,0,1,1,0,0,1,2,0,1,1,-1,1,-1,-1,-2,1,-1,-1,0,0,0,0,1,1,0,0,-1,-1,-1};
			448: counter1_out = '{0,-1,-1,2,-1,0,-1,1,0,2,-1,2,-1,0,-1,0,0,0,-1,1,0,-1,0,-1,0,1,0,0,0,2,1,-1,1,1,1,-1,0,-1,0,0,0,0,-1,1,0,-1,0,-2,0,1,-1,0,-1,-1,-1,-1,-1,0,-1,0,0,1,-2,-2,2,0,0,1,-1,0,0,1,1,2,-2,1,0,1,-1,0,1,0,-2,0,-1,0,0,1,-1,0,-2,1,0,-1,0,0,-1,-1,-1,2};
			449: counter1_out = '{-1,2,-2,1,0,1,-1,0,1,-1,0,0,1,1,0,0,-1,1,2,0,0,0,0,-1,0,0,-1,0,2,-1,-1,-2,1,1,2,0,-1,-1,1,1,2,0,-1,0,1,1,-1,0,-1,0,1,-1,0,-2,1,1,-1,1,-1,0,1,1,1,-1,-1,0,0,1,0,-2,-1,2,0,-2,0,0,-1,-1,0,0,0,0,0,1,0,-1,0,0,-2,0,1,-1,1,-1,0,1,2,0,0,1};
			450: counter1_out = '{-1,0,1,-1,0,0,0,-1,2,1,-1,3,0,0,-1,0,1,0,-1,-1,-1,1,-1,1,1,0,0,0,0,0,-1,1,2,1,0,0,-1,0,1,-1,0,-1,-1,1,-2,0,-1,-1,0,0,0,0,0,1,0,1,2,-2,-1,1,0,-1,-1,1,-1,1,-2,0,0,0,-1,-1,0,-1,-1,2,0,1,0,-1,1,1,0,0,1,-1,0,-1,2,0,0,1,-1,-1,-2,0,1,0,2,1};
			451: counter1_out = '{0,1,1,0,0,-3,-1,0,0,0,2,1,1,0,1,0,0,0,1,1,1,0,2,0,1,0,0,0,-2,1,-1,-2,0,0,0,-2,0,0,1,-1,1,-2,0,0,1,-1,1,1,-1,-1,0,-1,1,-2,-2,-1,0,1,1,1,-1,-1,-1,2,1,-1,-1,1,0,-1,-2,0,-1,-1,0,0,-1,0,-2,0,-1,1,-1,-1,-1,0,1,1,0,1,0,0,0,-2,-2,0,0,1,0,1};
			452: counter1_out = '{1,-2,1,0,-1,-2,1,1,1,1,1,-2,0,-1,0,-1,1,2,0,1,0,0,0,2,0,1,1,0,1,0,1,-2,-1,1,0,0,0,-2,0,-1,0,0,-1,0,-1,-1,0,0,-1,0,0,0,1,0,0,-2,1,0,-1,0,0,0,-1,0,1,0,-1,-2,0,1,1,0,0,0,-1,1,1,0,-1,-1,0,0,0,1,0,-1,0,1,0,0,0,0,1,-1,0,1,0,1,-2,-1};
			453: counter1_out = '{0,-1,0,0,-1,-1,0,1,1,0,1,0,0,-1,-2,0,0,0,-2,1,0,0,-1,1,0,0,0,-1,-1,0,-1,0,1,1,0,1,1,-1,0,0,1,1,2,-1,1,0,0,2,-1,-1,-1,-1,-1,0,1,0,1,-1,-1,0,2,0,-1,-1,-1,2,0,0,-1,1,2,1,-1,0,0,0,0,-1,1,0,2,0,-1,0,-3,0,0,0,0,1,-1,-1,1,1,1,1,1,1,-1,0};
			454: counter1_out = '{0,-1,1,0,0,1,0,-1,1,-1,0,-2,0,2,-1,0,1,-1,2,0,0,0,1,-1,0,0,-1,0,1,-1,-1,-1,1,0,0,-2,0,0,-2,-1,1,1,1,2,0,0,-2,0,-1,-2,-3,0,2,1,0,1,1,1,-2,2,-1,0,1,0,0,-2,-2,0,0,1,0,-2,0,1,-1,1,-2,0,-2,0,1,-1,-1,-1,-1,-1,0,0,-2,2,-1,-1,1,1,-2,-2,0,1,-2,-1};
			455: counter1_out = '{-1,1,3,1,0,0,0,-1,2,-1,0,1,0,0,1,0,0,1,1,3,1,0,0,0,-1,-2,1,1,1,1,-2,0,1,-1,0,-1,0,0,-1,2,1,-1,1,3,0,-2,-1,0,-1,-3,-1,0,1,-2,1,0,-1,-1,1,-1,1,0,1,1,0,1,-1,0,1,-2,1,0,2,3,1,1,-1,0,1,1,-1,1,-2,0,0,0,1,-1,0,-3,-1,0,-1,1,1,-1,0,2,0,-1};
			456: counter1_out = '{1,-1,0,-1,-1,1,1,0,0,0,0,-1,-2,1,1,-1,1,1,1,1,0,0,0,0,1,-1,1,0,-1,0,-2,0,-1,0,1,-2,0,0,0,0,-1,-1,0,1,-1,-2,2,-2,-2,-3,-1,-1,0,2,-1,0,-1,-1,1,-1,-2,1,2,0,0,-1,1,-2,0,-2,2,-2,0,0,-2,2,-2,1,-1,0,1,0,-1,3,-1,-1,-1,0,1,-2,0,-1,1,0,-1,1,0,0,2,0};
			457: counter1_out = '{0,-1,-1,0,0,1,0,-1,0,-1,1,1,0,-1,-1,1,-2,0,-1,-1,1,-2,1,0,0,-2,0,0,1,1,0,-1,0,1,-1,0,-1,0,0,-1,-3,0,0,1,2,1,0,1,-1,-2,-1,1,-2,-1,0,1,0,0,-1,-1,1,0,0,-1,2,-1,0,0,-1,-1,1,-1,0,0,1,0,-2,2,-1,1,1,0,-1,0,0,-1,0,0,1,-2,0,-2,-2,2,-1,0,-2,-2,0,0};
			458: counter1_out = '{0,2,1,0,-1,0,1,0,2,0,-1,-2,-1,0,1,0,0,2,0,0,0,1,0,0,0,1,0,1,2,3,0,-1,0,1,-2,1,1,-1,1,-2,-3,0,1,1,1,-1,-1,0,-2,-2,0,1,0,-1,-1,1,1,1,0,0,1,0,-1,0,2,-1,0,-2,0,-2,2,0,1,0,0,0,-2,1,0,-2,0,1,-2,1,-1,0,-1,-1,1,1,0,-1,1,1,-1,1,1,-1,0,0};
			459: counter1_out = '{3,0,0,-1,-1,0,-1,-2,-1,0,1,1,-1,0,0,-1,-1,0,1,2,-2,0,-1,0,-1,-2,-1,0,1,-1,0,1,-1,-2,1,0,0,-1,0,0,-1,2,-1,0,0,0,0,0,-1,-1,1,0,0,0,0,0,0,0,2,-1,0,0,-2,-1,-2,0,1,0,-1,-1,-2,0,0,-2,1,-1,-1,0,-1,-1,-1,-3,-1,-2,0,-1,0,0,1,1,0,2,-1,2,-3,0,-1,0,1,0};
			460: counter1_out = '{4,-1,1,-1,0,0,3,-3,0,1,1,1,1,1,2,-1,1,0,4,0,1,-1,1,-1,2,0,-2,-1,0,-1,2,0,0,1,0,0,2,1,0,-1,-1,3,-1,0,2,0,0,-1,-3,0,-2,-1,0,1,0,-1,-1,-1,0,0,-2,0,0,0,1,0,1,0,0,1,-1,-1,-1,-1,0,3,1,-1,-1,0,-2,-1,0,-1,0,-1,0,0,0,0,1,-2,-1,-1,-2,3,-1,0,2,1};
			461: counter1_out = '{0,-1,0,0,-2,-2,2,-2,2,0,-1,1,2,0,0,-1,0,-1,3,0,0,-1,-1,0,2,0,0,1,0,-1,1,1,0,0,3,0,-1,1,0,0,-2,1,0,2,1,0,-1,1,-2,0,-1,-2,0,1,0,0,2,-2,1,0,0,-2,1,0,0,2,0,2,0,-1,1,0,1,0,-1,0,1,1,-1,-1,-1,0,0,0,0,-1,0,1,1,0,1,-1,-1,-1,-1,1,0,0,1,-2};
			462: counter1_out = '{0,-3,2,0,0,-3,1,0,0,1,0,0,-1,1,-2,1,1,0,-1,0,-1,1,0,-2,1,0,-1,1,1,-2,2,0,0,-1,1,1,0,1,0,-1,-3,1,0,2,0,-1,0,0,-2,0,1,-3,0,0,2,0,2,-1,0,-1,1,-1,0,-1,0,-1,-1,-1,0,-1,1,1,1,0,0,-1,2,-1,1,1,0,0,0,-1,1,0,0,0,-1,1,-1,0,1,0,0,1,1,2,-1,-1};
			463: counter1_out = '{-1,-1,0,2,0,-1,-2,1,1,-1,0,0,-2,1,-1,0,0,0,0,1,2,3,0,0,2,0,0,0,0,-2,1,1,-2,0,0,-2,1,-1,-1,0,0,1,0,0,1,-2,1,0,-2,1,0,-2,-1,-1,0,1,0,-2,1,0,0,2,1,0,0,-1,1,-1,-1,-3,2,0,-2,1,-1,1,0,0,-1,-2,-3,0,0,0,1,-1,0,-1,1,-1,0,-3,-2,0,0,0,0,0,0,1};
			464: counter1_out = '{0,-1,2,1,0,0,1,0,-1,2,2,-1,-2,1,-1,-1,-1,1,-1,0,0,2,0,2,-2,0,-1,1,0,0,-1,-1,0,0,-1,0,-1,-1,0,1,-1,-1,0,1,1,0,2,1,0,1,1,-1,1,2,-1,2,0,0,1,0,-1,1,0,-1,1,-1,2,0,-1,1,1,-1,0,1,0,-1,0,-1,1,-1,0,1,-2,2,1,1,0,-1,2,0,0,-1,0,1,0,1,-1,1,-1,-1};
			465: counter1_out = '{0,2,0,-1,0,-3,1,0,0,-1,0,-1,-1,0,1,0,-1,0,0,1,1,1,0,2,0,-1,1,1,1,0,0,-1,1,-1,-1,-2,2,1,2,-1,-2,-1,-1,-1,0,-1,-1,-1,0,1,0,-1,0,-1,0,1,-2,-1,-1,-1,1,1,-2,0,-1,-3,2,-1,2,-1,-1,0,-1,1,1,0,-2,1,-1,1,0,-1,-2,0,1,0,-1,0,-2,-1,-1,-2,1,0,-1,-2,-2,1,0,2};
			466: counter1_out = '{1,-1,-1,0,-1,-1,0,0,0,0,0,0,1,-1,0,-1,1,-1,-1,1,1,0,1,1,0,0,1,0,0,-1,2,0,-1,0,0,-1,1,-1,0,0,1,-2,1,0,0,-1,0,-1,0,0,1,1,1,1,-1,1,-2,0,0,-2,1,0,0,1,0,2,0,1,0,0,0,0,0,2,1,2,-1,2,0,-1,-1,0,0,-1,-1,0,0,-1,-1,-2,0,-2,1,2,1,-1,-1,-1,0,-1};
			467: counter1_out = '{-2,-1,0,0,0,-2,-2,1,0,0,1,-1,0,1,0,-1,-1,0,-1,0,0,0,0,0,-2,-1,1,-2,2,1,0,-2,-1,0,0,0,0,0,1,0,-1,-2,1,-1,-1,-1,0,0,-2,0,-1,0,-2,0,-1,2,0,1,0,1,0,1,2,2,0,0,0,0,2,-1,0,-1,-1,2,1,2,0,2,1,0,-1,-1,0,-1,1,1,1,0,-1,0,0,1,1,2,-2,-2,0,-1,1,-1};
			468: counter1_out = '{-2,1,2,1,1,-1,0,1,0,0,-1,-2,2,1,-1,0,-1,0,0,-1,1,1,1,-1,0,0,0,-1,0,1,-1,-1,1,2,0,-2,1,-1,2,0,0,0,0,0,0,-2,-2,-2,0,1,-1,-1,1,-1,-1,0,1,-1,1,0,1,-1,0,1,0,1,0,-1,0,1,-1,-2,1,-1,1,0,-2,0,0,0,-3,-1,1,-1,2,-1,-1,2,-2,-1,-1,1,0,2,0,-1,-1,0,-1,0};
			469: counter1_out = '{0,-2,-1,-1,-2,-1,0,0,2,2,0,1,1,-2,1,0,1,0,-1,-1,0,-1,0,1,1,-1,1,0,0,3,1,-2,0,1,0,0,-1,1,0,-1,1,-2,0,-1,1,0,0,1,1,1,1,1,-1,0,-1,1,-1,0,0,-1,3,1,2,-1,0,0,-1,2,-1,1,0,0,-1,-1,0,3,0,1,-1,-2,-2,-1,0,0,0,0,1,0,-1,0,0,0,1,1,1,0,-1,0,0,0};
			470: counter1_out = '{-1,1,3,-2,1,0,-1,1,1,2,1,-1,1,0,0,0,0,0,0,0,-1,0,-3,0,-1,0,0,-1,1,-2,0,1,0,2,0,1,1,-1,0,0,0,1,-1,1,-1,-1,-2,0,1,1,-1,1,0,2,0,0,-2,0,-2,1,1,1,1,1,2,-2,0,-1,-1,0,-1,0,1,1,1,1,1,-1,1,-1,0,-1,1,0,0,2,-2,-2,0,-1,1,0,1,-1,-2,-2,1,-1,-1,0};
			471: counter1_out = '{1,0,0,0,-1,1,1,-1,-1,0,-1,0,0,1,-1,-2,-1,0,-1,2,1,-2,0,0,0,0,0,0,-2,0,1,0,0,0,0,1,0,1,1,-1,0,2,2,0,1,1,0,0,1,0,0,0,-1,-1,2,1,-1,-1,0,-1,1,1,1,0,3,-2,0,0,0,1,0,-1,-1,1,3,-1,-1,1,1,-2,-3,0,-1,1,0,0,1,1,-1,-2,-1,1,1,1,0,0,1,-1,0,2};
			472: counter1_out = '{0,0,1,-1,1,0,1,1,-1,0,0,0,0,0,0,0,0,-1,0,0,0,-1,0,-1,1,-1,-2,1,0,0,0,0,-2,-1,-2,-1,-2,0,0,0,-2,2,1,1,0,0,0,0,0,-2,-2,0,0,0,1,0,1,-1,-1,-1,2,0,1,0,1,0,-1,0,1,0,-1,0,1,-2,1,-1,0,0,-1,-1,-1,2,0,1,0,-2,2,-1,-1,0,1,-2,1,1,0,0,0,0,0,0};
			473: counter1_out = '{-1,2,1,1,0,0,2,0,1,1,2,0,0,1,0,0,-1,0,1,-1,1,-1,-1,0,1,0,-1,0,0,0,-1,-2,0,0,2,1,2,0,1,2,0,1,0,1,2,2,0,-1,-1,1,0,-1,-1,1,0,1,0,1,-1,1,-2,-1,0,-1,0,1,2,0,1,0,1,-1,0,-2,0,1,0,0,-1,1,0,-1,-1,-1,1,-1,-1,0,0,0,0,2,1,-1,0,-1,1,1,1,3};
			474: counter1_out = '{-1,0,0,0,2,1,0,-2,0,-1,-1,2,1,0,2,0,-1,-2,0,1,-1,0,-1,-2,-2,-1,1,-1,0,0,1,-1,1,1,0,-1,0,2,0,0,0,-1,0,0,0,1,-1,1,0,-2,0,-1,-1,0,1,-1,0,0,-2,0,1,1,1,1,0,-1,0,-1,0,0,-1,0,1,1,1,-1,0,0,0,0,-1,-2,-1,-1,-1,-1,1,-1,-1,-1,-1,-2,0,1,1,-1,-1,-1,-2,-2};
			475: counter1_out = '{1,-1,0,0,0,-1,-3,1,1,2,0,1,-2,2,-1,1,0,-1,2,0,1,1,-2,-1,1,-2,2,-1,0,-1,0,0,1,1,0,1,1,0,-1,1,-1,2,-1,0,1,0,0,0,0,-3,-1,0,0,0,0,1,-1,0,1,1,2,2,0,1,1,0,-1,2,0,1,0,0,0,-1,1,1,0,-1,-1,1,0,1,-1,2,0,2,1,-1,0,0,-1,0,1,-1,-1,1,0,-2,-1,0};
			476: counter1_out = '{0,1,-1,-3,2,0,-2,0,1,0,-1,1,1,0,-1,-1,-1,-2,1,-2,-1,1,0,-2,0,0,1,0,0,-1,-1,0,-1,0,0,2,0,-2,0,0,-1,1,-1,0,0,0,0,0,-1,0,-2,-1,2,0,0,0,1,0,1,0,0,0,-2,0,1,-1,-1,-1,0,-1,2,0,0,0,-1,0,2,0,2,0,0,0,-2,0,-1,1,-1,0,1,0,0,-1,0,1,0,0,1,2,1,0};
			477: counter1_out = '{0,-2,0,1,0,1,1,-1,1,2,-1,-2,0,0,0,0,0,-1,1,0,-1,2,-1,0,0,0,0,0,0,1,-1,0,-1,-1,0,-1,-2,-1,1,-1,1,0,-1,0,-1,-1,1,-1,0,-1,-1,-2,-2,0,-2,-1,0,-1,1,-2,-1,0,0,0,-1,1,-1,-2,1,-1,-1,-1,0,-1,0,1,1,1,-1,0,-1,0,-1,-2,0,0,0,0,0,-1,2,1,0,1,0,0,-1,-2,0,-1};
			478: counter1_out = '{0,-2,0,0,0,-1,-1,1,-1,0,1,-1,0,0,0,0,0,-2,0,-1,-1,1,1,-1,1,-1,0,1,-1,1,1,1,2,-1,1,2,0,0,-1,0,-1,0,1,1,1,2,-1,-1,1,2,1,1,0,1,0,0,1,1,-1,-1,-1,0,-1,1,0,1,0,-3,-1,0,0,0,0,1,1,-1,0,0,0,-1,0,0,-1,0,0,1,0,-1,-1,-1,-2,0,-1,1,0,1,0,1,2,0};
			479: counter1_out = '{0,1,0,0,0,1,0,-2,-2,3,-1,1,0,1,0,0,1,-1,0,1,-1,1,-1,0,1,1,1,-2,-1,-2,-1,1,-1,-1,-1,-1,1,2,0,0,0,-1,0,2,0,-1,-2,0,1,0,0,0,1,0,2,0,1,0,0,1,0,-3,-1,-1,0,-1,-1,-1,-2,-1,-3,0,0,-1,0,2,0,1,0,-1,-1,1,-2,0,-1,-1,0,-1,-1,-1,1,2,1,1,1,0,0,-1,0,1};
			480: counter1_out = '{1,0,-2,0,1,-1,1,-1,0,0,1,-1,0,-3,1,0,1,0,-1,1,-2,2,2,-1,0,-2,1,0,-1,-2,0,1,0,0,0,1,2,0,-1,1,1,0,0,0,0,-2,-2,0,0,1,1,1,0,-1,0,-1,0,-2,-2,-1,0,2,0,-1,0,2,-2,-2,0,-1,-2,-2,0,0,1,1,-1,-3,0,0,-2,0,1,0,0,0,-1,0,-1,-2,1,-1,0,-1,1,0,0,-2,-1,-1};
			481: counter1_out = '{1,1,-1,0,-1,2,-1,-1,1,1,0,0,1,0,1,-1,0,-2,1,2,0,-1,1,-3,-1,0,1,-1,-1,1,0,-1,0,-1,1,-1,0,0,0,2,0,-1,0,-1,0,0,-1,-1,0,0,1,2,1,-1,1,2,2,0,0,0,-1,1,-1,-1,1,0,-1,0,-2,2,-1,1,0,2,0,-1,-1,-1,0,1,1,-1,-1,-2,0,0,0,1,0,0,1,-2,2,0,1,1,1,0,-1,0};
			482: counter1_out = '{1,0,0,0,-1,-1,1,-1,-1,-1,0,0,0,0,0,0,1,0,-1,1,0,0,-1,1,0,1,1,1,-3,1,0,0,1,0,-2,1,-1,-1,-1,0,1,1,-1,2,1,-1,0,-2,0,-1,1,0,-1,0,0,1,1,2,-1,-1,1,0,1,-1,0,1,-1,-2,1,1,0,0,0,-1,0,3,1,-2,0,0,0,-1,1,0,0,0,0,0,-1,1,-1,-1,1,2,0,0,0,0,0,0};
			483: counter1_out = '{1,0,0,2,1,1,0,0,2,-2,0,-1,1,-2,-2,-2,1,-1,-1,1,-1,-1,0,3,-1,0,3,-1,-1,-1,-2,0,1,2,1,0,0,0,0,-1,1,-1,0,0,0,-2,0,-1,1,0,0,0,-1,0,2,2,0,-1,0,-1,0,1,-3,-1,1,-1,-1,1,0,0,0,-1,1,1,1,1,-3,1,-1,3,0,0,0,1,-2,0,-1,0,1,-1,-1,-1,0,1,-2,-1,-1,0,0,-1};
			484: counter1_out = '{0,1,1,-1,1,-1,-1,0,0,-1,-1,0,-1,-1,2,-1,-1,1,-2,1,-1,-2,0,0,-2,3,2,0,1,2,0,0,0,1,-1,-1,1,-2,-1,1,-2,-1,0,1,1,0,1,-1,-1,1,-1,-1,-1,1,2,0,0,0,0,0,1,-2,1,-1,0,1,0,-1,-1,-1,-1,0,0,2,0,0,-1,-1,0,2,-1,2,0,1,-1,1,0,0,2,-2,0,1,1,2,-1,0,-1,-1,2,1};
			485: counter1_out = '{0,-1,-1,0,1,0,0,-1,0,0,0,0,-1,0,-1,0,-1,0,1,0,0,0,-2,0,0,-1,-1,1,0,1,0,0,1,1,0,0,-1,0,0,-1,-1,-1,1,1,0,0,0,2,-1,-1,-1,-1,0,-2,1,1,1,-3,1,0,1,1,1,-1,1,0,-1,0,1,-4,0,-2,1,1,-1,-1,-3,0,0,-2,-1,0,0,0,-2,1,-1,0,-1,-2,2,0,0,1,0,0,0,2,2,-1};
			486: counter1_out = '{3,0,0,0,1,0,0,0,-1,-2,-1,1,0,-2,-1,-2,-2,-1,2,0,0,1,0,1,-2,-1,1,0,0,1,0,1,1,0,0,2,0,1,1,2,-2,-1,1,0,2,-1,0,-1,-4,-1,-1,-1,0,-1,1,0,2,0,1,0,0,0,1,0,-1,-1,1,0,1,-3,1,0,-1,-2,-2,0,-4,-1,-1,-3,3,-1,1,-1,-1,0,-1,-1,0,1,1,-2,-1,0,-3,0,1,0,3,0};
			487: counter1_out = '{2,-1,-2,-1,-1,0,1,-2,1,0,0,-1,-1,1,2,0,-1,-1,2,1,0,1,0,-1,0,0,-2,1,0,0,2,1,0,1,1,1,1,-1,0,-1,0,1,2,2,0,-1,0,0,-3,0,-1,0,-1,1,2,0,-1,1,1,0,1,1,1,1,1,-1,-1,-1,0,-2,2,1,-1,-2,-1,0,-2,1,-4,1,-1,0,-1,0,0,-3,0,0,1,1,2,-2,-1,2,-1,-1,0,2,-1,2};
			488: counter1_out = '{1,0,-1,1,0,1,-1,-2,1,-1,1,0,-1,1,2,-2,-2,-2,0,1,1,0,0,-1,0,2,-1,1,0,0,0,1,1,1,0,0,-1,1,0,-1,0,0,2,0,0,2,2,0,-2,-1,-1,1,1,-1,0,1,1,-1,1,1,1,-2,1,-1,1,0,0,-1,1,1,2,1,0,-1,1,0,-2,0,-3,0,0,2,0,0,-1,-1,0,1,1,1,2,-2,0,0,-2,1,-1,1,0,-1};
			489: counter1_out = '{1,-1,0,0,-2,0,1,0,1,1,1,0,-1,0,1,1,-1,-2,-2,0,2,1,0,-1,0,2,-2,0,1,1,3,-1,-1,0,0,-1,1,0,1,0,-1,3,0,1,1,0,0,1,-1,-1,0,-1,1,0,1,0,1,-1,0,-1,-1,-1,1,-2,2,0,-1,1,1,-1,-1,-1,0,0,-1,-1,-1,0,-2,2,0,-2,-2,1,-1,0,-1,1,2,1,-1,0,0,0,-2,-1,-2,-1,0,1};
			490: counter1_out = '{0,0,0,1,-1,-1,0,-1,0,-1,-1,-1,-2,0,0,0,1,-1,-1,1,-3,0,1,1,0,1,-1,1,0,-1,1,1,-2,2,-1,-1,0,0,1,0,0,2,-1,-2,2,0,3,-1,-3,-1,1,-1,0,0,0,2,1,-1,1,-1,1,-2,1,0,1,-2,0,0,-1,-2,1,0,0,3,1,1,-1,-2,-1,1,0,1,1,-2,-1,-1,-1,1,2,2,-1,-3,0,-1,0,-1,-2,1,1,0};
			491: counter1_out = '{0,1,1,1,2,0,1,-1,1,0,-1,0,-2,-1,-2,0,1,-1,0,1,0,1,0,3,1,-1,0,-2,2,1,0,-1,1,1,0,-4,1,2,-1,1,-1,0,0,2,1,1,-1,0,-2,1,0,-2,1,2,1,0,-1,-2,0,1,0,0,-1,-1,-1,0,0,0,2,-2,-1,1,1,1,0,0,-1,0,0,-2,0,1,0,-2,-1,0,-2,-1,-1,-1,-2,-2,-2,1,-1,-2,0,0,2,0};
			492: counter1_out = '{0,0,-1,0,-1,1,0,1,0,0,1,-2,0,0,0,2,-1,0,0,1,0,0,0,0,-1,0,2,2,1,2,0,-2,-1,-1,-1,-1,1,1,2,0,1,0,0,0,1,1,1,1,-2,-1,1,-1,0,1,1,1,-2,-1,0,0,0,0,1,1,1,-2,1,0,1,-1,0,-1,2,1,1,1,-2,1,-1,-1,0,2,-2,-1,0,0,0,1,0,1,0,0,0,-1,1,-2,1,-1,-1,0};
			493: counter1_out = '{0,0,-2,0,0,1,-2,-2,-1,1,0,1,0,-1,-1,1,1,0,-1,1,-1,-1,-1,0,0,1,2,-1,0,-1,0,1,0,-1,0,-1,-1,1,-1,-1,-1,-1,0,-1,0,-3,1,-1,0,-2,-1,0,3,0,0,0,-2,0,0,0,1,-1,-1,0,0,-1,-1,-1,4,-1,0,2,0,0,2,1,-1,0,0,-1,1,1,1,0,1,0,-1,-2,-4,0,-2,-1,-2,1,-2,-1,1,-1,0,-1};
			494: counter1_out = '{1,-1,-1,0,0,-2,0,-1,0,1,1,-3,1,0,1,-1,1,-1,0,0,1,-2,1,0,1,0,1,-2,0,-1,0,-1,0,1,0,-1,-1,0,1,0,-1,0,-1,-1,0,-1,0,1,-1,-1,0,1,2,3,-2,1,-2,2,-3,1,0,0,0,-1,-2,1,-2,0,1,-1,-1,1,-1,1,1,0,-1,0,0,-1,-1,2,-1,0,1,2,1,0,0,1,0,0,1,0,1,1,1,1,-1,-1};
			495: counter1_out = '{2,-2,-1,0,0,-2,1,1,1,2,-1,0,0,1,1,0,0,0,-1,0,-3,0,0,1,0,2,1,0,-1,0,0,-1,0,1,1,0,-1,0,2,-1,0,-1,0,0,-1,0,-2,1,2,1,0,0,-2,0,0,0,0,-1,-1,0,-1,0,-1,1,2,0,0,0,0,0,1,-1,1,-1,-2,1,-1,-1,0,1,1,-3,-1,2,1,1,1,0,-2,0,-2,-1,0,2,1,1,-1,-1,1,1};
			496: counter1_out = '{1,0,-2,-2,0,-2,1,1,0,1,1,0,-1,2,1,2,1,1,1,0,0,0,-2,0,0,1,0,0,-1,-1,-1,-1,1,0,-1,0,-1,0,-1,1,-1,-1,-1,1,-1,0,-1,-1,1,-1,0,2,-1,1,2,-2,0,2,-1,-1,0,0,0,-1,1,-1,0,0,2,1,2,0,0,1,1,0,0,0,0,0,-1,-2,-2,-2,0,-1,1,0,-2,0,-1,0,-1,0,0,-1,-1,1,1,1};
			497: counter1_out = '{0,-2,-1,0,1,0,1,-1,2,-1,1,0,1,0,0,0,0,1,1,1,-1,-1,1,1,1,1,1,1,-1,0,0,-1,-1,0,-2,1,0,-1,0,0,0,0,0,1,1,-3,0,-1,-1,-1,0,0,-2,0,-1,2,-1,-1,0,-1,-1,1,0,0,0,0,1,-1,2,2,1,1,1,0,1,0,-1,1,-1,1,0,-1,1,-1,1,-1,1,-1,0,1,1,0,-1,0,0,0,1,-1,-2,-1};
			498: counter1_out = '{-1,0,-1,-1,-1,1,0,0,-1,0,1,1,-1,1,-1,0,-2,1,2,-1,-2,1,0,1,1,-1,1,0,-1,1,0,-1,0,0,1,0,-2,-1,1,1,1,-2,0,-1,1,1,-1,1,1,-1,-1,0,1,-1,0,0,-1,1,-1,0,-1,0,1,-1,0,-3,0,-1,0,1,1,0,1,1,1,-1,1,1,-1,-1,-1,-2,0,-1,0,0,0,1,0,-1,1,1,3,0,0,-1,1,1,0,1};
			499: counter1_out = '{0,-2,1,2,0,0,0,0,-1,0,0,-1,0,1,0,1,0,-1,0,0,-2,0,-1,-3,1,-1,2,1,-2,-2,1,0,-1,-1,-1,3,0,0,-1,-2,-1,1,2,0,-1,0,-1,1,1,-1,-1,0,0,1,-2,1,-2,2,0,0,-1,0,0,-1,1,1,0,-1,1,0,1,-1,0,-1,2,-1,1,2,0,2,-1,-2,0,0,2,1,0,-1,-1,-1,2,-1,1,-1,-1,0,1,-1,0,-1};
			500: counter1_out = '{-1,0,-1,0,0,-2,1,0,-1,-2,-1,0,0,0,2,-1,0,2,2,0,0,0,0,1,0,-3,-1,2,-2,-1,0,0,0,-2,1,1,-1,-1,-1,0,-1,1,-1,0,-1,0,2,0,0,3,-1,0,0,-2,-1,1,0,0,0,-1,-1,1,0,1,-1,-1,0,0,-1,0,3,0,1,0,-1,1,1,-1,-2,0,-2,-2,1,1,0,0,3,0,-1,-1,0,-1,1,-2,-1,0,0,1,-1,0};
			501: counter1_out = '{0,0,1,0,0,1,-1,1,0,-1,-2,0,0,-1,0,1,2,-1,-1,-3,1,0,0,-1,-1,1,1,2,-2,0,0,1,1,-1,1,-1,1,1,-2,0,-1,1,-1,0,0,-1,1,-1,0,1,-2,1,0,1,2,0,-2,-1,-1,1,0,-2,0,0,0,-1,-1,-2,-2,1,0,1,-1,-2,1,-2,0,0,0,0,0,0,-1,-1,1,0,0,0,0,2,0,0,0,1,1,-1,0,-1,0,1};
			502: counter1_out = '{0,1,0,0,0,0,0,0,1,0,1,0,1,1,0,0,0,0,0,0,-1,0,1,1,0,-1,0,0,-1,-1,0,0,1,1,-2,-1,2,-1,1,2,1,-2,-2,1,1,0,1,0,0,1,-1,0,-2,-2,-1,0,1,-1,-1,2,2,-1,0,0,1,-1,0,1,2,-1,-1,-1,0,0,-2,0,-1,-1,-1,-1,3,-1,-1,0,0,2,1,-1,-1,0,0,1,1,1,1,0,0,-1,2,0};
			503: counter1_out = '{-2,-1,0,0,-2,1,2,-1,2,-1,-1,0,1,-2,1,1,0,0,0,-2,0,1,-1,-1,1,1,0,0,1,-1,0,0,0,0,0,0,0,0,0,1,0,1,1,-1,0,2,-2,1,0,1,2,-1,3,0,0,1,-1,-1,0,-1,1,0,1,0,-2,0,3,0,-1,-1,0,-1,0,-1,1,0,2,1,0,1,4,1,-1,-1,0,0,0,0,0,0,0,0,1,0,1,1,0,-1,1,-1};
			504: counter1_out = '{-2,2,-1,2,0,1,-1,0,-1,1,-1,-1,1,0,-1,-1,0,1,0,1,0,0,0,0,-1,1,0,0,-1,1,0,1,3,0,0,0,1,1,0,1,-1,-1,-1,-1,1,0,-2,-1,0,1,-1,1,-2,1,0,-1,0,-1,0,0,0,0,-1,-1,-2,0,-1,0,0,-1,0,0,0,1,1,-1,2,-1,0,1,0,1,3,-2,-2,-1,0,-2,-1,-1,0,0,-1,1,0,1,1,1,2,-1};
			505: counter1_out = '{-1,-1,0,-1,0,0,0,-1,0,-1,-1,0,-2,1,0,1,1,2,-1,-1,0,-1,-1,0,-2,1,-1,1,1,0,-1,-1,1,-1,1,1,2,-1,-1,0,0,-1,1,1,0,-1,0,-1,0,-1,0,0,0,0,0,-1,2,1,0,1,0,0,2,0,-1,1,1,0,-1,0,1,1,0,1,0,0,-1,1,0,2,-1,-1,-1,0,-1,-1,0,1,1,-1,1,2,1,-1,0,-1,0,0,0,1};
			506: counter1_out = '{1,1,-1,2,0,0,0,1,0,1,-2,-1,-1,0,-1,-2,1,-2,0,-2,1,0,1,0,1,1,0,1,0,1,1,-1,0,2,-1,-1,-1,0,-1,0,0,1,-1,2,-1,1,0,0,-1,2,0,-1,1,-1,0,0,1,0,0,0,-2,0,0,0,-1,0,0,-1,0,1,0,0,2,0,0,0,1,1,1,1,-2,-1,0,2,0,-1,0,-1,0,2,-1,-1,2,0,1,1,0,0,-1,0};
			507: counter1_out = '{-1,-1,1,-1,1,-1,2,-1,1,0,0,0,-1,0,0,-1,0,0,-1,0,-2,0,0,1,1,-1,0,1,-1,-1,0,1,1,0,0,-1,-2,0,1,1,1,-1,0,-2,1,-1,0,2,1,-2,0,1,-2,1,-2,1,0,1,1,0,-1,1,0,1,0,1,3,1,-2,2,0,-1,-3,0,0,-1,0,-2,0,1,-1,-1,0,0,0,0,2,0,-1,1,2,1,0,0,0,-1,1,-1,-2,0};
			508: counter1_out = '{0,-1,-3,0,0,-1,0,0,0,1,0,2,0,0,0,0,2,0,0,0,-2,1,0,1,-1,1,2,0,-2,1,0,0,2,0,2,-1,2,-1,1,0,-1,-2,0,0,-1,0,1,0,-1,1,2,1,0,-1,0,-1,1,1,2,0,1,-1,0,1,0,-1,0,-2,2,0,2,-1,0,-1,1,-1,-1,-1,0,0,-1,0,1,0,-1,-2,0,-1,-1,-1,1,2,-1,1,0,-2,2,0,-1,0};
			509: counter1_out = '{2,1,-1,2,-1,-1,-3,-1,0,-1,0,0,1,0,0,1,-2,0,2,1,0,1,0,2,0,1,2,0,-1,-2,1,-1,0,-1,1,2,-1,-2,1,-1,0,1,1,-1,0,-2,0,0,-1,-1,-2,0,1,1,-1,0,-1,-1,-1,-1,2,1,-1,1,0,-1,0,-1,1,2,1,-1,1,-1,2,1,1,0,0,-1,-1,-1,-1,0,0,-1,3,-1,1,-2,1,-2,0,0,1,0,0,0,-2,1};
			510: counter1_out = '{2,0,0,0,0,-2,1,1,1,0,0,1,1,-1,-1,-1,0,0,1,2,-1,0,0,1,-1,0,1,-2,0,0,1,1,1,2,0,-3,-1,0,0,2,1,2,0,-1,0,1,0,0,0,0,-1,1,0,-1,1,0,1,-1,0,0,-1,-1,0,1,0,0,0,-1,-1,-1,-1,-1,1,1,0,1,2,-1,0,-1,-1,0,-1,0,-1,-1,-1,-1,-1,1,-1,-1,2,0,0,-1,0,2,0,0};
			511: counter1_out = '{0,1,-1,1,2,-1,0,0,-1,-2,1,0,-1,0,0,-2,1,-1,-2,1,-2,0,0,0,-2,-2,2,-1,-3,0,-1,1,3,1,-1,-1,-1,0,0,-1,3,-1,1,1,1,-1,0,0,0,-1,-1,1,-1,-1,0,1,-2,-1,0,1,1,0,-1,-2,1,0,0,-1,-1,-2,-1,0,0,0,1,2,-1,0,-1,0,1,-2,1,2,0,0,0,-1,1,0,-2,-1,-1,-1,-2,-1,0,2,0,1};
			512: counter1_out = '{2,-1,0,-1,0,1,-2,-1,-1,-2,1,0,0,0,0,-2,3,0,1,0,1,0,0,1,-1,-1,1,-2,-2,1,-1,1,0,-1,1,-2,-1,0,-2,0,1,-1,0,-1,0,0,-1,0,1,0,-2,1,0,0,1,0,0,0,-1,1,0,1,0,1,2,1,1,0,0,-1,-1,2,-1,1,1,-1,-1,-1,-1,0,1,1,-1,-1,-2,-1,0,0,1,1,1,0,1,1,-1,-1,1,-1,2,1};
			513: counter1_out = '{3,2,-1,-1,0,-3,1,0,0,-2,-1,0,0,-2,0,-1,1,0,1,2,1,0,-1,0,-2,0,0,1,-2,4,0,0,-1,0,1,0,0,-1,1,0,4,-1,0,0,1,-1,2,0,-2,0,-2,1,0,1,-1,-1,0,-1,0,-1,1,0,0,0,-1,1,1,-1,1,-1,-1,0,0,-2,1,-1,-1,0,0,0,-1,-1,-1,0,-2,-1,-1,-1,0,-1,-1,0,-3,1,-1,-1,0,1,1,0};
			514: counter1_out = '{2,2,-1,0,1,0,0,-2,-1,-1,1,-1,0,1,0,1,0,-1,2,0,1,-1,-1,-1,-3,-1,0,-1,-2,1,-1,0,0,-1,2,1,-2,-1,1,-2,1,-1,2,0,1,0,1,1,0,0,-1,0,0,1,1,2,-1,-1,1,0,2,-2,1,0,0,0,1,0,0,-1,1,1,-1,-1,1,0,0,-3,-1,0,0,0,-1,0,-2,-1,1,-2,0,1,0,1,1,1,-1,0,-1,-1,0,1};
			515: counter1_out = '{2,0,1,1,0,0,1,-1,0,-2,0,0,0,-1,1,1,0,2,1,0,0,2,-1,-3,-1,1,0,1,0,0,1,1,0,0,1,0,0,-1,0,-2,-2,-1,-1,0,2,0,1,0,1,-3,-2,-1,1,0,-1,-1,0,0,2,1,1,0,0,0,1,0,-1,1,1,-1,0,1,-2,-1,-1,-1,-1,-1,0,-1,-1,0,1,1,-2,-3,-1,-2,0,-1,-1,1,-2,-1,-1,-2,-2,-1,1,-1};
			516: counter1_out = '{0,-1,0,0,1,-1,2,-2,0,0,2,1,-2,1,0,0,-1,-1,0,0,-1,1,-1,-3,-2,0,-1,1,0,-2,0,-1,-3,-1,0,0,0,-1,2,0,1,2,-1,2,1,-2,0,-1,-1,-1,-1,-4,-2,-1,-1,-1,0,-1,0,0,0,1,0,1,0,0,1,0,0,-1,-1,0,-1,-1,1,-1,-2,-1,-2,0,0,0,0,-2,-2,-1,0,-1,2,1,2,-1,-1,0,0,-2,-1,0,1,0};
			517: counter1_out = '{0,-1,0,1,2,-1,1,-2,0,0,2,-1,-2,1,2,-1,-1,-2,-1,1,1,-1,1,0,-1,0,0,0,-2,0,1,-2,1,-1,0,-2,-1,-1,1,1,0,2,-1,0,-1,0,1,1,-1,-2,-2,-1,0,0,1,1,0,1,0,0,0,-1,0,-1,0,-1,-1,0,-1,-1,0,1,2,0,1,-2,-1,1,-1,0,-1,-1,-2,1,-1,3,0,0,2,1,-1,0,-1,-2,1,1,1,-2,2,0};
			518: counter1_out = '{0,0,-1,0,2,-2,1,1,-2,-1,0,-1,-3,1,0,1,-1,-1,-1,-1,-2,-2,-2,3,0,1,2,0,-2,-1,-2,-1,1,1,0,-2,-1,-1,-2,1,1,0,1,2,0,0,-1,-1,-2,0,1,-1,0,4,2,1,-1,1,0,0,0,-1,0,1,1,0,3,0,2,0,1,0,2,1,1,-1,0,-1,-1,-2,-1,-2,0,-1,0,0,-2,0,0,0,-3,-1,1,-1,-2,-2,-1,0,0,0};
			519: counter1_out = '{-2,0,1,0,1,-1,-1,0,-1,1,0,-4,-1,-2,1,0,1,0,1,0,0,-2,0,-1,-1,-1,2,1,-2,-2,0,-2,1,0,0,-1,-1,0,0,1,-1,0,-1,1,-1,-2,1,1,-1,0,1,-1,0,3,-1,0,-1,0,-2,0,-1,-3,-1,-1,-1,-2,1,2,0,2,0,0,0,1,1,-1,-1,0,-1,1,0,0,2,0,0,0,-1,2,-4,0,0,0,-1,1,-1,0,-1,1,0,0};
			520: counter1_out = '{1,2,-1,2,-2,-1,0,-1,1,0,-1,-2,2,1,0,-1,-1,0,1,0,1,-1,1,0,0,1,1,0,-1,1,-2,-1,1,0,-1,-3,-1,-1,0,0,1,0,0,0,-1,0,-2,0,-2,-1,-1,0,1,1,-1,0,-3,1,1,0,1,0,-1,0,-1,-3,-1,-2,1,-1,-2,1,1,0,1,1,0,2,1,-1,-1,-1,1,0,0,0,-1,0,0,-1,-2,-2,0,2,-1,-2,-2,-1,-1,0};
			521: counter1_out = '{-1,0,1,2,1,0,-2,1,1,0,-1,-2,1,-1,1,0,-1,-1,-2,1,0,0,0,2,-1,0,0,-4,-2,0,-1,-2,2,-1,0,0,1,1,1,2,1,0,1,1,1,0,-2,1,-1,1,1,0,1,0,-1,0,-1,0,-1,-1,-1,0,-1,-1,1,1,0,1,0,-1,0,0,1,-1,1,1,0,1,0,-1,-1,2,1,0,1,1,1,-1,0,1,-1,-1,1,1,0,-2,2,0,0,1};
			522: counter1_out = '{1,1,-2,0,0,-1,-1,0,1,2,0,1,1,0,0,0,0,0,-2,1,-1,0,0,0,-1,-2,0,-1,-1,1,1,-2,0,-1,0,0,0,0,1,0,-2,-2,0,-1,1,0,0,0,0,0,1,0,-1,-2,1,0,-3,-1,0,0,-1,1,2,1,0,1,2,-1,1,0,0,2,-1,1,0,-1,-1,2,0,0,-3,0,0,0,0,0,-1,1,0,-1,0,-1,1,2,-1,0,0,1,-1,0};
			523: counter1_out = '{-1,1,-1,0,0,-1,1,-1,1,-1,1,-1,-1,2,-1,-1,-3,-2,0,1,0,0,0,-1,-1,1,-1,1,-2,-1,-2,0,0,1,0,1,-2,0,1,1,1,-1,0,1,0,2,-1,0,0,1,1,-1,-1,-1,-1,0,-1,1,-2,0,1,2,0,-2,1,2,0,0,0,1,-2,2,-1,-1,-1,1,-1,0,0,0,-1,0,0,-1,0,-1,1,1,0,0,-1,-1,0,1,-1,-1,-1,-1,-1,-1};
			524: counter1_out = '{1,-1,1,0,1,0,-1,0,0,1,0,0,0,-1,-1,1,0,1,2,0,0,0,1,-1,0,-1,-1,-1,-1,0,-1,1,-1,1,1,1,1,0,0,1,-2,-1,-2,-1,-1,0,-1,-1,1,1,0,1,-1,0,1,2,0,1,0,-1,0,1,-1,0,1,-3,0,0,1,0,0,1,-1,-1,0,-1,0,1,0,0,-2,0,-1,1,1,0,-1,0,-1,0,-1,0,-2,1,0,2,1,1,1,1};
			525: counter1_out = '{0,-2,-1,-1,1,0,0,2,1,0,1,-1,-1,0,1,1,0,0,-1,3,1,-1,-1,-1,0,0,2,-1,1,-1,1,0,-3,1,1,1,1,0,1,-1,1,-3,-2,0,0,-1,1,0,1,1,-2,-2,-2,0,0,-2,-2,1,1,0,0,1,0,2,-1,0,1,0,1,1,0,0,1,2,1,-3,0,0,0,-1,-1,-2,-2,-1,0,-1,1,0,1,0,0,1,-1,-1,1,0,1,1,-3,-1};
			526: counter1_out = '{0,-1,1,-1,1,0,0,-2,1,2,0,0,1,1,-2,1,0,0,0,-1,-1,0,1,0,0,0,0,1,0,1,-1,-1,0,0,1,1,0,0,0,0,0,-1,-2,0,1,1,0,0,1,2,1,1,1,-1,0,0,-2,0,0,1,0,1,-1,1,-3,0,0,-1,0,2,2,0,0,0,0,0,-3,0,-1,1,1,-1,1,2,0,-2,0,-1,1,0,2,1,2,1,-3,-1,1,-1,1,-1};
			527: counter1_out = '{-1,2,0,0,0,0,1,0,0,-1,1,1,1,-2,-2,-1,0,-1,1,-1,-2,1,-3,0,1,-3,-1,0,-1,0,0,-1,2,1,1,0,-1,-1,1,0,0,1,0,1,0,-1,-1,0,-1,0,-2,-1,-2,-1,0,1,-1,-2,0,0,0,-1,-1,0,2,-1,-1,0,1,1,0,0,-1,0,2,-2,1,0,0,0,0,0,0,0,-2,0,0,-2,1,-2,1,-1,0,-1,0,-1,1,-2,1,0};
			528: counter1_out = '{0,1,1,-1,-1,1,-1,0,-1,-1,0,0,0,-1,2,0,1,1,2,0,-2,0,1,2,1,1,0,1,0,-1,-2,-2,-1,2,-1,0,2,1,1,0,0,-2,0,1,-2,1,2,-1,0,1,-1,0,-1,0,2,0,0,1,1,1,-2,0,0,0,3,-1,1,0,0,-3,-2,-1,1,-1,0,0,0,-2,0,0,0,1,0,0,-1,-1,3,0,2,-1,1,0,2,0,0,0,0,0,-1,-1};
			529: counter1_out = '{0,-2,0,1,0,-1,2,1,-2,0,0,-3,-1,0,1,1,1,-1,0,-1,0,2,0,0,1,-1,0,0,-2,0,-2,1,0,-1,1,1,0,0,0,1,1,0,-1,1,0,0,2,0,0,1,0,-2,-1,1,0,0,0,-1,-2,1,-1,1,1,-1,0,0,-1,-1,0,0,-1,1,0,1,0,-1,0,-1,2,0,-1,-2,1,0,0,1,-1,0,1,0,0,-1,1,-2,0,0,0,-1,0,1};
			530: counter1_out = '{0,0,0,0,1,-2,-1,-1,0,-1,0,0,-1,0,1,0,2,1,0,1,1,0,2,-2,-1,0,-1,0,-2,-1,0,0,-1,0,0,-1,-1,1,0,0,-1,0,0,1,1,-2,-2,2,-1,-1,0,-1,0,0,1,-1,1,0,0,-1,2,-1,1,0,1,-1,0,0,1,-1,0,-1,0,-3,-1,0,2,0,-1,0,0,0,1,0,-3,0,-1,0,-1,-1,-1,1,-1,0,-2,1,2,1,0,0};
			531: counter1_out = '{-1,0,0,1,2,1,-2,1,1,1,1,1,0,-1,1,-1,1,0,1,-1,2,0,0,0,0,0,0,0,-1,1,1,-1,0,-1,-1,2,1,-1,-2,2,0,1,-1,0,1,1,0,1,1,0,-1,-1,-1,0,-1,1,1,0,1,0,0,0,-1,0,0,0,0,0,1,1,0,0,-1,0,-1,0,0,0,-1,-2,0,-1,0,1,-1,-1,0,0,0,1,1,1,0,-1,0,-2,0,2,-2,1};
			532: counter1_out = '{1,1,0,-1,0,-2,1,0,0,0,-1,0,0,-1,-3,-1,-2,0,-1,1,0,1,-1,0,0,1,-1,-1,0,0,1,0,1,0,0,0,-1,1,0,-1,2,1,0,-1,-1,0,1,-1,2,0,-1,0,0,0,1,-1,0,-1,0,0,0,-1,1,-2,-1,0,-1,-1,1,2,1,1,1,1,0,1,0,-1,-1,0,0,1,-1,0,-1,0,2,-1,0,-1,-2,0,-1,-1,-1,-1,0,-2,1,0};
			533: counter1_out = '{0,0,0,-2,-1,0,0,0,0,0,1,1,0,2,0,1,0,0,-1,0,-2,0,1,2,-2,-1,1,0,2,0,-1,-1,0,0,-1,1,0,0,0,0,0,0,-2,0,-1,-1,-1,0,-1,-1,0,-1,0,-2,1,2,-2,0,2,0,1,1,-1,-1,1,0,-2,2,2,1,0,1,0,2,1,0,0,-2,2,0,0,1,-1,0,-1,-1,1,-1,0,-1,3,-1,0,0,0,0,2,1,-1,1};
			534: counter1_out = '{1,1,-1,1,-1,-1,0,-1,-1,0,-2,1,-1,0,2,0,0,0,-2,1,-1,0,0,0,-2,0,-1,1,0,0,1,2,0,-1,1,0,0,-1,0,3,1,0,0,0,0,0,1,0,0,0,-1,0,-2,0,0,0,0,-1,1,-1,1,-1,0,1,1,0,0,0,1,0,-1,-1,-1,1,2,-1,0,-2,-2,-1,0,-2,0,1,-1,-1,0,1,-1,1,1,0,1,0,-1,0,0,-1,-1,1};
			535: counter1_out = '{3,2,0,2,-2,-1,-2,-1,0,2,0,0,0,0,-1,-2,0,1,0,0,0,-1,0,0,0,-1,0,1,1,-1,0,0,1,-1,0,1,0,-1,1,0,1,0,2,1,1,-2,-1,2,0,2,0,-1,-2,1,-2,2,-2,0,-2,0,-1,1,-1,0,0,-1,0,2,3,1,0,-1,-1,0,2,-1,1,1,2,1,1,-1,-2,1,1,0,0,0,-1,1,-1,1,1,-1,1,2,0,0,0,-1};
			536: counter1_out = '{1,1,0,0,0,1,0,1,1,-1,1,1,0,1,1,-1,-2,1,0,0,2,0,1,0,1,1,0,1,-1,1,0,-1,1,-1,0,-2,2,0,-1,2,1,-2,1,2,-1,1,0,-2,0,1,0,0,1,1,0,1,0,0,0,-1,2,1,-1,-1,-2,1,-1,0,-1,1,-2,-1,0,0,1,2,0,1,0,-2,0,0,0,-1,2,0,1,0,0,0,2,2,-2,1,-2,0,1,1,-1,-1};
			537: counter1_out = '{0,-1,-1,0,1,-1,2,0,-1,1,1,0,0,0,2,-2,0,2,-1,2,0,-1,1,0,0,-1,1,0,-3,1,-1,-1,1,0,-1,1,-1,0,-1,2,1,0,-1,0,1,-3,-1,0,1,2,1,0,1,1,1,0,-1,-1,0,0,0,2,0,-1,0,0,1,0,1,2,1,1,-1,1,0,1,0,0,0,1,0,0,1,0,-1,-1,2,0,0,0,-1,2,1,1,-1,-1,1,0,0,-1};
			538: counter1_out = '{1,0,0,0,-1,-2,1,1,0,-1,-1,1,0,1,0,-2,0,-1,-2,1,-1,-2,0,1,0,0,1,0,-4,2,1,-1,1,0,1,-2,-1,2,0,-1,-1,-2,-1,1,0,-2,1,-1,1,3,-1,0,0,-2,0,1,0,-1,0,-1,-1,-1,0,1,1,1,1,-3,1,1,1,-1,-1,0,1,-1,2,0,0,0,-2,1,-1,-1,-1,0,0,-1,0,0,-1,1,-1,-2,-2,0,-1,-2,-1,1};
			539: counter1_out = '{2,-1,1,1,1,0,-1,-1,-1,1,1,-1,-1,2,0,0,1,1,0,0,0,0,0,-2,-1,-2,2,0,-1,2,0,-1,0,0,1,-2,-2,0,0,0,1,-1,0,-1,0,0,1,1,-1,2,-1,-1,0,1,1,1,-1,-1,-1,-2,-2,1,-2,-1,-1,1,1,-1,0,2,0,0,1,0,0,1,-2,0,1,2,-1,1,0,-1,0,-1,1,0,1,-1,0,0,2,0,-1,-1,1,0,1,1};
			540: counter1_out = '{3,0,-2,0,0,2,0,0,-2,-1,0,1,-1,1,0,0,1,-1,1,0,-1,0,1,0,-2,-2,0,0,-6,2,-1,1,1,-1,-1,0,0,1,0,0,1,1,3,0,0,2,1,-2,0,0,0,1,1,0,1,0,1,0,0,-1,1,1,0,-1,-1,0,1,1,0,-2,0,0,-2,0,2,0,1,-2,0,0,0,-1,-1,-1,0,-2,1,0,0,1,2,-1,0,0,-1,0,0,1,0,1};
			541: counter1_out = '{2,1,0,-1,0,-1,0,1,1,1,0,-1,1,0,0,0,-2,0,2,1,-1,-2,0,1,-2,0,-1,2,-4,2,-2,0,0,1,1,0,0,-1,-1,0,0,1,0,1,1,-1,1,2,1,0,-1,0,0,1,0,0,0,2,-2,-1,-2,-1,1,1,-1,0,0,1,1,-2,0,-1,0,0,-1,-2,0,0,1,2,0,1,0,-2,1,-2,0,0,1,-2,0,0,1,1,-1,2,1,0,-1,0};
			542: counter1_out = '{-1,-2,-1,1,0,-2,0,0,0,0,2,1,0,0,2,-1,1,0,3,-1,1,-1,-1,-4,-3,0,-2,2,-7,-1,-1,1,0,-1,1,1,-2,0,2,0,1,0,0,0,2,-1,0,0,0,0,-1,-1,0,1,0,1,1,-2,-3,0,-1,1,1,-1,0,-1,1,1,-1,0,-1,-1,-1,-3,0,-1,0,1,0,0,1,-1,1,-1,-1,0,-2,-1,0,0,-1,-2,0,1,0,0,1,1,-1,1};
			543: counter1_out = '{0,1,1,0,1,-1,1,-3,-2,0,2,0,2,0,1,0,0,-1,0,-1,0,0,0,-2,-4,1,1,1,-4,-2,0,0,1,0,0,1,0,0,1,0,1,-2,0,-1,0,-1,2,0,-1,1,-1,0,-1,2,1,-2,1,1,-1,1,1,1,-1,0,1,-1,1,2,2,0,0,1,-1,-3,1,0,-2,0,-1,1,0,-1,0,1,-1,0,-2,-1,0,1,1,0,-1,3,-1,1,0,1,1,1};
			544: counter1_out = '{1,1,-1,-1,0,1,3,-1,-1,0,-1,1,-1,0,2,0,0,0,0,0,1,2,0,-3,-2,3,1,1,-3,-1,0,0,0,0,-2,0,1,0,0,1,1,-1,0,3,-1,1,1,0,0,-1,-1,-1,2,-1,2,1,2,0,-1,0,2,1,-1,0,0,1,0,-1,1,0,0,1,-1,0,1,-1,-1,1,-1,-2,0,0,0,-2,-1,1,-1,0,2,1,1,1,0,0,0,-1,0,0,0,1};
			545: counter1_out = '{0,2,1,1,1,-1,1,-2,-3,-1,-1,0,-1,0,0,0,-1,-1,-2,-1,1,0,1,2,-2,1,-1,2,-2,-1,1,0,1,0,-1,-2,1,0,-1,0,3,-1,2,1,0,1,-1,-1,0,1,-3,0,1,0,2,1,2,-1,-1,-2,1,0,0,-1,0,2,1,0,-2,-2,-1,-2,1,1,1,-1,1,1,1,-1,0,0,2,0,-1,-1,-1,1,1,2,0,1,0,-1,1,0,0,1,0,1};
			546: counter1_out = '{-1,2,-1,0,0,1,2,-1,-2,-3,-1,0,-2,-1,0,-1,0,-1,-1,-3,0,-1,0,2,0,0,0,1,-1,0,1,0,0,3,-1,0,-1,0,-1,-2,2,-1,1,0,-1,1,0,1,1,0,1,-1,2,4,0,-1,0,-2,-1,1,0,-1,-1,-1,0,-2,-1,-1,0,0,0,0,1,0,0,1,-2,-1,-1,0,-1,0,0,0,2,-2,0,-1,-2,0,-2,1,1,0,1,1,0,1,1,1};
			547: counter1_out = '{1,0,-1,2,-1,0,-1,1,-2,-1,0,-1,0,0,1,-2,-1,-1,0,0,-2,-2,1,3,0,0,0,1,-1,-2,0,0,-1,1,1,2,0,0,0,-2,0,1,0,0,-1,0,0,0,-1,2,-2,0,2,3,1,0,-1,-2,0,1,0,1,0,0,0,-2,1,-2,2,1,0,1,0,1,1,0,0,3,0,-1,1,-1,0,-1,1,-2,0,0,-2,-1,0,-1,1,-1,-1,-2,1,0,1,1};
			548: counter1_out = '{0,1,1,1,0,0,0,1,-1,-1,-2,-2,1,1,-2,1,0,-1,0,0,0,0,0,1,1,-1,0,1,0,0,0,-1,0,1,1,2,1,0,0,1,1,1,0,1,2,-2,0,0,1,-1,-1,0,2,0,0,-1,-2,1,-2,0,-1,-1,2,0,1,0,1,-1,0,1,-2,0,1,-1,1,1,-1,1,-1,-2,0,-1,0,1,2,-1,-1,0,-2,-1,-1,-1,-1,1,0,0,0,0,-1,-1};
			549: counter1_out = '{-1,1,0,1,-1,3,-1,0,1,-1,0,0,-1,1,-1,-1,2,-1,2,-1,1,-2,0,1,0,1,0,1,-2,0,0,0,0,-1,0,2,-1,-1,1,0,-2,-1,-1,-1,-1,-2,0,-1,0,2,1,0,0,-2,-1,0,0,0,0,-1,0,-1,-2,-1,-1,0,0,-1,1,3,1,3,-1,-1,1,1,-2,-1,-1,0,-2,-3,0,1,-1,1,0,0,-1,1,-2,-2,-1,-2,1,0,-1,2,0,1};
			550: counter1_out = '{1,-2,-1,0,2,-2,0,-1,0,1,0,2,0,0,1,0,-1,0,0,2,-2,0,0,-1,-1,0,1,1,0,1,0,3,-1,1,1,0,-2,1,-1,1,0,3,1,1,1,2,1,1,0,-1,-1,0,0,0,-2,0,-1,-2,-2,3,1,2,-1,-1,0,2,-2,-1,1,3,0,1,1,0,2,1,-1,1,1,-2,-1,0,-1,0,-1,0,1,1,-1,0,-1,2,-1,0,1,-3,1,1,0,1};
			551: counter1_out = '{1,-2,-1,-2,0,-2,-2,1,2,0,2,0,0,0,-2,1,-1,-1,-1,1,0,-1,0,0,0,1,-1,1,-1,-2,-1,-1,0,1,0,2,1,0,0,2,0,-1,0,-1,1,2,0,0,0,0,-1,-1,-1,0,-2,0,-1,0,-2,2,0,0,0,-1,2,0,1,2,2,-1,0,1,-1,-2,-1,0,0,0,0,0,-2,0,-1,2,0,-1,-1,-2,1,2,-1,0,0,-1,1,0,0,0,2,0};
			552: counter1_out = '{0,-1,1,0,-1,0,-1,-1,1,0,-1,0,0,-1,0,1,-2,2,-2,0,1,-2,0,-1,1,0,1,1,0,0,0,1,2,1,0,0,-1,-2,-1,1,-1,0,-1,0,1,2,1,1,-1,1,-1,2,-1,0,0,1,0,0,0,1,-1,1,0,1,3,2,1,1,0,0,0,0,0,-1,-1,-1,0,1,-2,0,0,1,1,2,1,0,-1,-4,0,0,0,0,-1,1,1,-2,1,0,0,0};
			553: counter1_out = '{0,-1,-1,-2,-1,-1,0,-1,2,0,1,2,-1,-1,0,-1,0,-1,1,-2,0,0,-1,-1,0,1,0,2,-1,0,2,1,-1,0,0,-1,-1,0,0,-1,-1,0,1,1,0,-1,1,0,1,1,-2,0,-1,0,0,0,-2,1,1,2,0,-1,0,-1,0,-1,-1,-1,1,-3,1,1,0,-1,1,-1,-2,0,-1,0,0,0,-1,0,0,-2,0,1,-1,-2,2,-1,2,0,0,0,1,-1,-1,0};
			554: counter1_out = '{0,-1,0,-1,1,0,-1,1,1,2,0,0,-2,2,-1,2,1,1,-2,0,-1,1,0,0,0,1,2,-1,0,0,3,-2,-1,0,1,0,-1,-1,0,-1,0,-1,-1,0,2,-2,-1,1,1,2,0,1,1,0,0,-2,-1,0,-2,-1,-1,1,0,-2,1,-3,0,-1,-1,-1,1,1,-2,-2,0,0,0,2,-1,-1,1,2,1,0,-2,-1,-1,-1,1,-1,1,-1,2,1,0,0,2,-1,1,1};
			555: counter1_out = '{-1,-1,-1,1,-1,-1,-2,-1,-1,0,-2,0,1,0,2,2,1,1,1,-1,-2,-1,2,0,0,-1,1,0,1,0,0,0,2,0,-1,0,0,1,0,0,1,0,0,0,3,-1,-2,1,-1,-1,-2,0,-3,1,1,1,1,-1,-1,0,-3,-3,-1,-2,1,0,0,-2,-1,0,2,0,-1,1,1,0,0,0,1,1,0,0,-1,-1,-2,0,-1,0,1,0,0,0,1,0,0,0,1,1,1,-2};
			556: counter1_out = '{2,-1,-1,2,1,1,-2,-1,-2,-1,1,-2,-1,-2,0,-1,0,-1,1,0,1,0,0,2,-1,1,0,1,0,-1,2,-2,1,0,-2,2,2,0,-1,-1,0,2,0,1,2,0,0,0,-1,0,0,0,-2,1,0,1,-1,0,0,0,-1,-1,0,-1,0,0,-1,-1,0,1,3,0,-1,0,0,-2,1,0,2,-1,0,-1,-1,-3,-1,1,1,1,0,0,-2,0,0,1,0,0,1,0,-2,0};
			557: counter1_out = '{0,0,-1,0,0,0,0,1,0,-1,0,0,-1,0,-1,0,2,1,0,0,0,2,1,-1,0,-1,0,-1,0,1,-1,1,0,1,1,1,0,-2,2,0,1,0,-1,-1,2,0,0,2,0,0,0,1,-3,2,1,0,2,-1,1,-2,0,0,-2,1,0,0,-1,2,0,0,1,0,0,1,0,-2,1,0,1,-1,0,0,0,1,1,1,-1,-1,0,0,1,1,1,-1,0,-1,2,-1,-1,0};
			558: counter1_out = '{1,1,2,1,1,0,0,0,-1,0,1,1,0,0,2,2,0,0,1,3,-1,0,0,2,2,0,-1,0,0,0,1,1,-1,1,-1,-1,-1,-2,1,0,-1,1,1,0,-1,0,2,1,-1,-1,0,0,0,1,-1,1,1,-2,1,-2,0,1,-1,-1,2,1,0,-2,-1,0,-1,1,1,0,0,0,1,2,2,0,1,0,0,0,0,1,0,1,4,0,1,-1,-1,0,-1,-1,0,1,-1,2};
			559: counter1_out = '{0,-1,1,0,0,0,0,0,0,1,1,-1,0,1,1,1,0,-1,-1,-1,0,1,1,1,2,1,0,0,1,0,-1,1,0,0,2,-2,2,-1,0,-1,-1,0,1,2,0,1,-1,1,1,0,0,0,-1,0,1,0,0,-1,1,0,1,1,1,-1,0,0,-1,1,0,0,-1,0,0,2,-1,1,2,-1,1,0,-1,0,1,0,0,-1,1,0,1,-1,-1,-1,0,-1,0,-2,1,0,0,-1};
			560: counter1_out = '{-2,0,0,0,0,-2,-1,1,0,2,-1,1,-1,1,-1,0,0,1,1,0,2,1,0,-1,0,1,1,1,1,1,0,1,2,0,-1,-2,-2,0,0,2,1,-1,1,1,1,0,1,-1,-1,0,1,-1,0,0,1,0,-3,1,-1,1,2,0,0,0,2,0,0,1,0,0,-1,1,0,-2,-1,0,1,-1,1,-1,1,-1,1,1,0,0,0,0,-1,0,0,1,1,1,-2,0,0,0,0,1};
			561: counter1_out = '{1,2,0,1,1,2,1,1,0,-1,0,2,0,1,1,-2,-2,-1,1,1,0,-2,2,1,-1,0,-1,0,-1,-3,0,-1,1,0,2,0,0,0,0,0,0,-1,0,0,1,-1,0,1,0,0,1,1,0,0,0,1,1,0,0,-1,-1,0,1,0,0,-1,-1,0,-1,1,1,-1,1,0,1,0,-1,1,0,0,-1,0,1,1,-2,0,0,1,0,0,-1,1,1,0,1,1,1,0,1,-1};
			562: counter1_out = '{0,1,1,0,0,1,-1,0,-1,1,1,1,1,-1,0,1,0,0,-1,-2,-1,-1,2,-1,1,-1,0,0,0,0,1,-1,1,0,3,2,0,1,-1,0,-1,0,-1,-1,0,-3,0,-1,1,-1,2,2,-1,2,1,-1,-1,-1,0,-2,-1,0,0,0,0,0,-1,1,1,-2,1,1,0,-1,0,-1,0,0,0,0,-2,0,2,-1,2,0,-1,-1,-1,0,0,0,1,0,1,1,0,-1,-1,0};
			563: counter1_out = '{1,-1,0,1,0,-1,1,1,1,-1,0,0,0,0,-1,1,0,1,1,-1,0,0,0,-1,0,0,1,0,1,-1,2,0,1,1,2,0,0,1,1,2,-2,-1,0,1,0,2,-1,-1,0,0,1,0,0,0,2,-1,1,1,-1,-1,0,-1,-1,-1,0,1,0,-1,0,1,1,0,1,-1,2,1,1,0,-1,-1,2,2,1,0,0,1,0,2,1,1,0,1,-1,-1,1,1,1,0,-1,0};
			564: counter1_out = '{3,-1,0,-1,-2,1,-2,1,0,-1,2,-2,-1,0,-1,-1,-2,0,-1,1,-2,1,1,-2,1,-1,1,1,-1,-1,1,1,2,-1,0,0,0,0,1,0,0,-1,1,0,0,1,0,0,0,-1,-2,-1,0,2,1,1,0,0,-1,0,1,0,0,-1,2,1,0,-2,-2,1,0,-2,0,-2,2,-1,2,2,0,1,0,0,1,1,1,-2,0,0,1,0,-1,1,0,0,1,1,0,-2,-1,0};
			565: counter1_out = '{0,1,0,-1,1,0,2,0,-1,-2,-1,0,-1,1,1,1,1,0,-1,-1,0,-1,1,-1,1,1,0,0,-3,0,-2,1,1,1,-2,0,0,2,-3,1,1,-2,1,0,1,-1,1,1,1,2,0,-1,2,-2,-2,-1,0,0,-1,1,-1,1,1,2,1,0,1,0,1,1,-1,0,1,0,0,1,0,0,-2,0,0,-1,1,0,1,0,1,0,0,-2,1,-2,0,1,1,-1,2,0,-2,1};
			566: counter1_out = '{2,1,-2,0,0,-1,1,0,0,0,1,0,0,-1,-2,0,-1,-1,0,-2,0,-1,-1,0,0,0,0,0,-2,1,-1,-1,1,0,1,-1,-2,1,-1,0,0,0,-1,1,1,-2,-1,1,0,3,1,0,1,-1,-1,0,0,-1,0,0,-1,-1,-1,-2,-1,2,1,-1,1,-2,-1,-1,1,-1,1,1,1,-1,1,1,-2,-1,0,0,1,-2,0,0,1,1,-2,2,-1,1,-5,0,-1,1,1,1};
			567: counter1_out = '{1,1,-2,1,0,-2,0,0,0,-2,-1,-1,-2,0,1,0,0,-1,1,0,0,0,-1,1,0,0,0,1,-3,3,1,1,1,-1,0,0,0,1,2,-1,0,-1,0,1,-1,0,0,0,1,1,0,0,0,0,0,-1,1,1,-1,-2,0,-1,0,0,-2,0,-1,-1,-1,1,-1,-2,1,1,1,1,3,-2,2,0,-1,1,-1,1,1,-3,0,0,0,-1,1,0,1,0,1,0,1,2,-1,-1};
			568: counter1_out = '{0,0,-1,0,1,0,3,1,-1,0,0,-1,2,0,1,0,2,0,1,0,0,1,0,1,0,1,0,0,-4,1,1,2,2,-1,1,0,0,1,-1,-1,-1,0,1,0,0,-3,1,0,2,2,-2,-1,0,2,0,1,3,-1,-1,0,0,0,0,1,-1,-1,0,0,0,1,2,2,0,0,3,1,1,2,1,0,-1,-1,1,-1,-1,0,-1,0,0,0,0,0,-1,0,0,0,0,-1,1,0};
			569: counter1_out = '{0,0,0,1,3,0,-1,0,0,0,0,1,1,-1,0,-1,0,0,2,0,-2,0,0,0,1,-1,1,-1,-3,2,1,1,0,-1,0,0,0,-1,2,2,1,-3,-1,2,-1,0,1,0,1,1,-1,0,-1,-1,0,-1,0,-1,0,0,-1,0,-2,2,-1,0,-1,1,0,1,-1,0,-1,-3,0,-1,0,3,0,0,1,-1,0,0,1,-1,1,0,-2,0,0,0,-1,-1,1,-1,-1,2,0,2};
			570: counter1_out = '{0,-1,0,-1,2,1,0,-1,0,0,0,0,-2,-2,-1,-2,-2,-2,1,-3,0,-3,0,-2,-1,0,1,1,-2,-1,1,0,2,-1,-1,-1,-2,1,0,-2,0,0,1,-2,0,0,1,0,-1,1,-2,-1,1,-1,1,0,0,0,0,0,1,0,-2,1,1,0,-1,0,1,0,2,0,-1,0,1,-1,1,1,1,-1,1,0,3,-2,0,-2,-1,1,1,1,0,1,2,0,0,0,1,-1,-2,-1};
			571: counter1_out = '{1,0,0,-1,1,-1,1,0,-3,0,1,0,1,2,0,-2,0,1,0,0,-1,-2,2,-2,-2,1,0,0,-3,0,-1,-1,1,2,0,1,-2,0,2,0,1,-1,2,1,1,-2,2,0,1,1,0,0,0,0,1,-1,1,-1,-1,1,-1,-1,-1,0,0,2,-1,-2,0,-2,1,1,-1,-2,0,-1,-1,3,1,0,2,-1,2,-1,1,0,0,-1,1,-1,-1,1,1,1,0,1,-1,-1,-1,0};
			572: counter1_out = '{0,-2,0,0,1,-2,2,0,-1,0,-1,0,-1,1,1,0,-1,0,1,-2,2,-1,0,-2,-3,2,0,2,-2,-1,2,1,2,1,0,1,0,0,1,-4,0,0,2,1,1,1,0,1,0,2,-1,-1,-1,1,1,0,1,0,0,1,0,1,-1,1,0,1,0,0,-2,2,-1,-1,0,1,-1,-1,-2,0,3,2,1,-1,2,0,-1,0,-1,-1,2,1,-1,2,0,0,0,4,1,0,0,1};
			573: counter1_out = '{-1,1,-3,1,1,1,1,0,-2,-1,-1,1,-1,-1,0,-1,-2,1,-1,-1,0,-1,0,1,0,0,0,2,-2,-1,1,0,0,2,-1,2,-1,1,1,1,1,-1,0,1,-2,-1,1,0,-1,0,-1,1,-2,0,0,-1,-1,-1,0,-1,0,2,0,0,0,-2,-1,1,1,2,-1,-1,0,-1,-1,-2,0,0,0,0,1,1,0,-1,1,0,-1,-1,0,0,0,1,1,0,0,0,2,-1,0,1};
			574: counter1_out = '{1,-2,0,1,2,-1,0,-1,-3,0,0,0,-1,1,0,-1,0,-1,-1,0,0,-2,1,3,1,0,2,2,-1,0,0,0,1,0,1,1,1,2,1,0,1,0,1,-1,0,-1,0,-2,0,0,-1,0,0,1,-1,0,0,0,0,0,1,1,-1,-2,0,0,-1,-2,-1,1,0,0,0,2,0,1,0,0,0,0,0,-2,0,1,0,0,0,1,0,-1,-1,-2,1,1,1,0,0,-1,0,0};
			575: counter1_out = '{0,0,1,1,1,0,-1,-1,-1,0,-1,0,1,0,-1,-1,2,2,0,1,0,0,0,1,0,0,1,0,-1,-2,1,0,2,0,1,2,1,1,2,-1,0,1,0,1,1,-1,1,-1,0,0,-2,-1,0,1,1,-2,1,2,0,1,-1,-1,0,0,-1,1,1,1,0,-1,-1,2,1,2,-1,0,0,1,-2,-1,-1,0,-1,1,1,0,1,1,0,1,0,-2,1,0,0,1,0,0,1,2};
			576: counter1_out = '{0,-1,1,1,0,0,0,-1,1,-1,-1,0,1,1,0,0,-2,-1,-1,-1,-2,-2,-1,1,-1,2,1,2,0,0,0,0,1,0,2,3,0,-1,-1,-1,-1,1,3,-2,2,-2,0,1,0,1,0,1,-1,-1,0,-1,-1,1,-1,0,2,1,0,-1,-1,0,1,0,0,-1,-1,-1,0,-1,-3,0,-1,1,1,-1,1,0,0,1,-1,-1,0,0,1,0,-1,-1,0,-2,0,0,0,0,-1,0};
			577: counter1_out = '{-1,0,0,2,1,2,0,0,0,-1,0,1,0,1,0,0,0,1,0,-1,-2,-1,1,0,1,0,0,2,-1,-1,2,1,1,-1,-1,1,0,0,0,2,0,-1,0,1,2,-2,1,-1,0,1,-1,0,-1,2,-1,-1,-1,0,1,-1,-1,-1,1,0,1,-1,1,2,0,0,-3,2,1,0,1,0,1,2,1,1,-1,1,1,0,0,1,0,1,-1,0,1,0,1,0,0,1,2,0,1,-1};
			578: counter1_out = '{0,-1,0,-2,0,1,0,0,2,0,-2,-2,-1,-1,-1,0,1,1,0,1,2,-1,0,-1,0,2,1,0,0,1,0,2,2,0,-2,1,-2,-2,-1,0,0,1,1,1,0,0,1,0,0,2,0,-1,-2,0,0,1,0,0,-1,1,-1,1,-1,-1,0,-1,-2,0,0,1,-1,0,0,0,2,-1,-1,-1,-1,0,0,-1,0,0,1,-2,2,1,-1,0,-1,1,1,-1,0,-1,3,0,1,0};
			579: counter1_out = '{-2,0,-1,-2,1,-1,1,0,0,0,1,0,0,1,-1,-1,0,1,0,0,-1,1,1,1,-1,0,1,0,-1,-1,0,1,1,1,1,1,1,0,1,1,0,0,0,-1,0,0,3,-2,0,0,1,-1,-1,-1,2,0,-1,0,0,-1,1,-2,-1,1,0,-1,1,1,0,0,-1,-1,-1,0,0,-2,-2,2,0,0,-1,0,-1,1,-1,-1,1,0,0,0,2,-2,1,0,-2,0,1,1,1,0};
			580: counter1_out = '{0,-2,-1,1,0,1,-1,0,2,1,-1,1,0,0,0,-1,0,0,-1,0,-1,-2,1,0,0,0,0,0,-1,-1,2,1,-2,1,3,0,-1,-1,1,1,-1,-1,0,0,1,-1,1,0,0,1,1,0,-2,2,0,0,-2,1,-1,-1,-1,0,1,1,1,-1,0,0,-1,-2,0,1,-3,-1,0,0,0,1,0,1,1,0,-1,0,-1,-2,0,0,1,-2,1,-1,-1,-2,-3,-1,1,0,-1,0};
			581: counter1_out = '{1,0,0,1,1,-1,0,1,-1,0,-2,1,0,0,1,1,0,0,-3,1,1,0,1,-2,1,-1,1,-1,1,-2,0,-2,0,-1,2,1,1,-2,0,0,-1,1,0,0,0,-1,0,0,0,2,0,0,-1,0,0,2,2,0,-1,1,-1,1,0,-1,2,0,-1,2,0,1,1,-1,-1,0,0,0,0,0,1,-2,-2,-1,-1,1,0,-2,0,-2,-1,0,0,0,1,-1,-1,1,1,1,-1,1};
			582: counter1_out = '{1,-1,0,0,0,-1,0,-1,0,1,-1,1,1,1,1,-1,1,-1,-1,-1,-2,-2,0,-1,-1,0,2,2,1,1,-2,0,0,-1,-1,0,-1,1,1,-1,-1,1,1,2,0,-1,1,0,0,0,-2,-1,0,1,-1,0,-1,1,-1,0,0,-1,1,0,1,-3,1,-2,0,0,1,0,-1,-1,1,-1,1,-1,0,0,1,1,0,-1,0,-2,-1,-1,0,-2,2,0,1,-1,-1,0,0,-1,0,1};
			583: counter1_out = '{-2,-1,-2,-1,0,0,0,-1,0,2,2,0,-2,-2,0,1,0,-1,2,0,1,2,1,0,-2,1,0,0,-1,1,0,0,1,-1,0,0,0,-1,1,-1,1,-1,1,2,0,2,1,0,0,3,-3,-2,-2,-1,1,-1,-1,2,0,1,0,2,-2,1,0,0,1,-1,1,1,2,1,0,-1,0,0,-2,0,0,0,0,0,0,-2,0,-1,-1,-1,-1,0,0,1,1,1,-1,-1,2,-2,2,0};
			584: counter1_out = '{0,1,-1,1,0,0,-2,0,0,0,-1,0,1,-1,-2,-1,1,2,1,1,0,0,0,2,0,0,2,0,0,1,-1,1,1,1,0,0,0,-1,1,1,1,1,0,0,1,-2,1,0,-1,-1,-1,-1,1,1,-1,0,1,0,0,1,1,-1,1,1,-1,1,-1,0,0,-1,-1,-1,-1,-1,2,0,-1,-1,2,-1,-1,1,1,1,0,0,1,-1,0,1,-1,0,-1,-3,0,1,1,-1,-2,1};
			585: counter1_out = '{0,0,2,-1,0,1,1,-1,0,1,-1,0,1,0,0,0,1,-1,1,1,1,-1,2,-1,-1,0,1,0,0,1,2,0,1,-2,0,1,0,0,0,0,-1,0,0,0,1,0,-1,0,0,-1,2,0,1,-3,1,-1,0,1,-1,1,-1,-1,0,-1,-1,1,-1,1,0,-2,1,2,1,-1,1,-2,2,-2,1,3,2,-2,-1,-1,0,0,0,0,-1,0,1,-1,0,0,0,0,0,-1,-1,1};
			586: counter1_out = '{0,1,0,0,-1,0,-1,-1,0,2,0,0,0,-1,0,-1,2,0,2,-1,1,1,0,2,-2,-1,1,0,1,1,-1,0,-1,0,0,0,2,0,-1,0,0,1,0,-1,0,0,0,0,1,1,2,0,0,-1,1,-1,0,1,1,1,2,0,1,0,0,-1,-2,0,-1,0,1,-1,-1,0,1,-2,0,-2,-1,1,0,-2,-2,-1,0,0,-1,0,1,-1,0,0,-1,0,0,0,3,2,0,-2};
			587: counter1_out = '{0,-2,1,1,1,0,-1,-2,0,0,-1,-1,0,1,1,0,-1,0,1,0,0,1,0,-2,-2,1,1,-2,-1,0,1,1,-2,1,0,0,2,-2,-1,0,1,0,-2,1,-1,0,0,-1,0,0,-1,-1,-2,-1,-1,0,1,0,1,-2,0,0,2,-2,-1,1,0,2,-1,-2,-1,-1,1,0,1,0,1,1,0,0,-2,-2,-1,2,-1,0,0,0,0,1,0,-1,-2,1,0,0,-1,-1,-1,1};
			588: counter1_out = '{-1,1,1,-1,1,1,0,-1,-1,0,0,-1,-1,-2,-1,-1,1,1,0,0,0,0,0,1,0,1,-1,0,-2,0,0,-1,-1,1,1,-1,2,1,0,-1,0,-1,1,0,-1,1,1,-1,2,1,2,0,-1,0,-1,1,0,-1,-1,1,-1,0,-1,-1,0,0,1,0,-1,0,0,2,1,-1,0,2,-1,-1,0,0,-1,1,0,0,-1,0,1,1,-1,-1,-1,-1,1,2,-2,1,1,0,1,1};
			589: counter1_out = '{0,0,-1,1,2,1,0,0,0,-1,0,2,2,1,2,-1,0,0,0,0,1,-1,1,0,-1,1,0,-1,1,1,1,1,1,0,-1,1,0,0,-1,0,0,1,1,1,-3,-1,0,0,0,-1,-1,0,1,0,0,-2,0,0,0,-1,0,1,-1,2,2,-2,-1,1,3,0,-2,0,0,0,-1,0,0,-1,1,1,0,0,0,1,0,-1,-1,-1,-1,-1,0,1,2,-1,0,0,0,0,-1,1};
			590: counter1_out = '{0,2,0,2,1,-1,0,0,2,-1,0,-1,0,2,-2,0,2,-1,1,0,0,2,0,-1,2,-1,0,1,1,-3,-2,-2,1,0,0,0,0,1,-1,0,0,1,-1,0,2,0,0,0,1,0,1,-1,1,0,-1,0,0,0,0,1,-1,0,-1,1,-2,-1,-1,0,0,-2,0,1,-1,0,-1,1,1,0,2,-1,-1,-1,1,1,0,0,-1,0,-1,0,0,-1,1,0,-1,0,-2,0,0,1};
			591: counter1_out = '{1,-2,1,0,1,1,0,2,1,1,1,2,1,1,-1,0,1,-1,1,0,-1,0,0,1,0,0,1,1,1,2,0,0,1,0,1,-1,2,-1,0,0,1,1,-1,1,0,0,0,1,0,-1,1,0,-1,0,1,1,0,0,0,0,-2,-1,-2,1,-1,0,2,0,1,0,-1,0,-1,0,0,0,0,-1,-1,-1,3,1,0,-1,0,0,1,-3,0,-1,0,2,1,1,-2,2,0,0,0,1};
			592: counter1_out = '{1,-1,-1,1,-1,-1,0,-1,1,0,1,-1,-2,1,1,1,1,-1,0,-1,-1,-1,1,0,2,1,2,0,1,0,-1,-2,0,0,-1,0,1,-1,-1,-1,-2,1,0,0,-1,-1,0,1,-1,3,0,0,0,0,-1,2,0,-1,-1,-1,-1,0,2,1,0,1,1,-1,2,0,1,1,-2,1,1,1,0,-2,0,0,1,-1,0,0,1,1,0,0,1,0,0,0,-1,-1,-1,-1,1,0,-1,-1};
			593: counter1_out = '{0,1,-2,0,0,0,0,0,-2,0,-1,0,-1,1,0,0,0,-1,1,-1,0,-2,0,-1,0,1,0,-2,0,1,0,0,0,-1,-1,0,1,-1,0,0,-1,0,1,0,1,0,0,-1,0,3,-1,1,1,-1,1,-1,-2,1,-1,-1,-1,1,-2,0,-1,0,-1,0,1,0,0,-1,1,0,-1,3,1,0,3,0,0,0,1,3,-1,0,0,-1,1,0,1,-1,0,0,-1,-2,1,1,-2,-1};
			594: counter1_out = '{0,-1,-1,0,0,0,0,2,1,1,1,0,0,-1,0,-1,0,-1,1,1,0,-2,-1,0,0,0,-1,0,-2,0,0,0,1,-3,0,2,0,0,0,1,0,0,-1,0,0,-1,0,-1,0,0,2,0,0,-1,1,-1,1,0,-2,1,-1,1,1,0,-1,0,1,2,1,1,-1,1,1,1,-1,0,-1,1,-1,0,1,0,0,-2,1,-2,0,0,0,1,0,1,0,0,-2,0,0,-1,0,1};
			595: counter1_out = '{1,2,-2,1,0,0,2,0,0,0,1,0,0,0,0,0,0,1,2,-3,0,-3,1,0,1,0,0,0,-1,2,0,-1,0,1,2,-1,2,1,0,0,0,-1,1,-2,1,-1,-1,1,-1,1,0,-1,0,0,1,-1,2,-2,-1,0,-2,0,-1,-1,-2,1,0,0,2,2,-2,-1,1,0,0,0,-1,1,1,0,1,0,1,0,-1,-2,0,-2,0,0,0,-2,-1,-2,2,0,-1,0,-2,0};
			596: counter1_out = '{0,-1,-2,2,0,0,-1,3,-1,1,1,-1,1,-1,-1,-1,0,-1,0,-1,-2,-2,0,1,0,1,1,-1,2,1,0,1,1,1,0,0,-1,2,0,-1,-1,2,1,1,0,0,0,1,-1,2,0,-1,-1,1,1,1,0,0,-1,-1,-1,1,-1,-1,1,1,0,1,1,0,0,-2,-1,-1,0,0,0,0,2,1,-1,2,1,1,0,0,-1,0,1,0,0,1,0,0,-1,0,0,1,1,0};
			597: counter1_out = '{0,2,0,-2,-2,0,0,1,-2,0,1,2,-1,-1,0,-1,0,-1,0,1,-1,-3,0,-1,2,-1,0,-1,1,0,0,-1,3,1,0,-1,-1,1,0,0,0,0,0,-1,0,0,1,0,-1,-1,0,-1,0,2,-1,0,0,1,-1,-2,0,1,0,2,0,1,1,1,0,2,0,1,-1,-1,0,0,0,1,3,2,-2,1,0,1,-1,1,-2,1,3,-2,0,0,-1,1,-2,-1,0,-1,-1,-1};
			598: counter1_out = '{-1,1,0,0,1,0,1,3,-1,-2,0,-1,1,1,-3,0,1,0,0,0,-2,0,0,0,0,0,-1,0,2,2,1,2,2,1,0,1,0,-1,0,1,-2,0,3,0,0,-1,0,0,1,2,1,-1,0,1,1,0,1,1,0,-3,-1,-1,1,0,-3,0,1,0,2,0,0,-2,-1,0,1,1,0,0,1,0,0,0,1,-1,-1,1,1,-2,0,0,2,-1,-1,1,0,1,0,0,-1,2};
			599: counter1_out = '{0,0,0,1,1,3,1,1,-1,0,1,0,-1,-1,1,-1,-2,-1,1,1,1,-1,0,-4,1,1,1,-1,1,-2,1,1,0,1,-2,0,0,1,0,1,2,-1,-1,0,-2,-2,1,0,-2,2,-1,1,1,3,0,-1,2,0,-3,-1,0,1,0,1,0,-1,0,-2,0,1,0,-1,-1,1,-1,1,-1,-1,2,2,0,-3,0,-1,0,0,2,-1,1,1,0,0,0,0,2,0,-2,1,0,0};
			600: counter1_out = '{1,0,1,0,1,0,2,1,-2,1,0,-1,-3,0,0,0,-2,0,1,-1,1,0,-1,-1,0,0,1,0,0,-2,1,-1,1,-1,0,-2,0,1,0,0,0,-1,2,1,0,0,0,1,0,1,0,-1,-1,2,-2,-2,0,-2,-1,-2,2,2,-1,1,-1,-1,2,-2,0,0,1,0,-1,0,1,-3,-1,0,-1,0,0,-2,0,-1,0,0,0,1,0,-1,0,-1,-2,1,1,-1,1,-1,0,0};
			601: counter1_out = '{-1,1,1,1,-1,1,0,0,0,0,0,-1,1,0,0,-1,0,-1,0,0,0,-2,-1,1,1,0,0,1,-1,-1,1,2,2,0,-1,0,1,-1,2,-1,0,-1,2,0,1,-1,1,1,-1,1,-1,0,-1,0,-2,-2,0,-2,-1,0,0,0,0,-1,-1,0,2,-1,1,1,0,0,0,0,0,0,-1,2,0,-1,0,-2,1,1,1,-2,2,0,-1,-1,1,0,0,0,-2,0,1,0,0,0};
			602: counter1_out = '{2,0,-1,0,-1,3,-1,1,-2,-1,0,2,1,-2,-1,-2,-1,0,-1,0,-2,-2,0,-2,0,1,-1,-2,0,0,-2,-1,0,0,1,2,-1,0,1,0,1,-1,1,-1,0,-1,0,1,1,0,0,0,2,0,0,-1,0,0,0,-1,-2,1,-1,-2,1,0,-1,-1,1,0,-1,0,1,1,0,-2,2,0,-2,-1,0,-1,0,2,1,-3,2,-2,-2,0,1,-2,-1,0,0,1,0,-1,0,2};
			603: counter1_out = '{0,-1,-3,0,1,0,1,0,1,1,0,1,0,0,0,0,1,-1,-1,0,-2,-1,0,2,2,1,1,1,0,-2,1,0,0,-1,1,1,0,2,1,-1,0,0,2,1,1,1,-1,0,2,1,1,-2,1,-1,-3,-2,2,2,-1,-2,0,1,-1,-2,0,0,-1,-1,0,1,-1,-2,0,-1,-1,0,0,0,0,0,1,1,1,-1,0,0,1,0,0,0,0,1,-2,-1,0,1,0,-1,0,0};
			604: counter1_out = '{0,1,0,2,-2,0,0,-1,0,0,-1,2,-1,-2,-1,-1,1,-1,0,0,-2,0,-1,1,-1,-1,-1,1,0,0,0,-1,0,2,1,0,0,0,0,0,0,-1,0,-1,0,1,1,-1,0,0,1,1,0,-1,-2,1,-1,0,0,-1,-1,1,-1,0,-2,1,-1,-2,0,1,1,-1,0,1,0,-1,0,-1,-3,1,0,0,2,-2,-1,2,0,0,-2,0,-1,0,0,-1,-1,1,-1,-1,0,-1};
			605: counter1_out = '{-1,-2,-2,-1,0,1,-1,0,0,-3,0,0,2,-1,-1,1,2,1,0,-1,-2,0,2,0,2,0,0,1,0,1,-1,1,1,-2,1,1,1,1,-1,1,-1,1,-1,0,0,0,1,-1,-1,1,0,1,0,1,-1,-2,1,0,-1,0,1,0,0,-2,1,-1,3,0,-1,-1,0,0,2,-2,-1,1,0,1,-1,-1,0,-2,-1,1,0,0,-2,-3,1,0,3,-1,0,-1,-1,1,1,1,-1,2};
			606: counter1_out = '{0,-2,2,0,0,0,-2,0,0,0,0,1,-1,1,0,1,0,1,1,0,-1,-1,-1,-1,1,0,-1,0,-1,1,0,0,0,1,1,1,2,-1,2,0,-1,1,1,1,1,-1,1,1,0,0,-2,0,-3,-2,0,1,-1,0,-1,0,0,0,2,0,-1,-1,0,0,1,1,0,2,0,1,-1,-2,0,1,0,1,-1,2,2,1,1,-1,-2,1,0,-1,0,0,0,0,-2,2,-1,-1,0,0};
			607: counter1_out = '{0,-1,-1,0,0,-1,-1,-1,0,1,0,-1,-1,-2,0,1,1,1,-1,-2,0,1,1,1,0,2,1,0,-1,1,-1,0,1,0,1,2,0,1,1,0,-2,0,-1,-1,0,0,0,0,0,1,-1,0,-2,2,1,-1,1,0,-1,0,-2,-1,1,-1,1,2,1,1,0,1,-1,1,-1,-1,1,0,-1,0,0,-1,-1,1,-1,0,0,0,0,-1,-2,-1,0,1,0,-2,0,-1,1,0,-1,-1};
			608: counter1_out = '{0,-2,-2,-2,0,1,-1,0,-1,-1,2,0,0,-1,0,0,3,-1,-1,1,0,1,1,1,2,1,2,0,0,0,1,-1,1,0,0,1,0,-1,0,0,2,0,0,-1,1,0,0,0,0,0,-2,1,0,-1,-1,2,-2,-1,-1,1,-1,-1,-1,1,3,0,-1,0,0,0,1,1,1,0,0,1,0,-1,2,-3,2,0,-1,2,1,-1,1,0,-2,0,1,1,1,-1,-2,1,1,-2,-2,-1};
			609: counter1_out = '{2,0,0,0,0,0,0,1,1,0,0,-3,0,0,1,-2,2,0,0,0,0,0,1,0,-1,0,1,1,-1,2,1,-1,1,-2,0,1,0,1,-2,0,-1,0,1,2,2,1,1,0,-1,1,0,0,1,-1,2,-1,1,0,-1,-1,-1,-1,0,-1,0,1,1,1,0,1,0,0,-1,0,-1,1,-1,0,-1,1,-1,1,-2,-2,1,-2,2,1,1,-1,-1,-1,1,0,0,1,1,0,-2,1};
			610: counter1_out = '{-1,-1,1,0,0,-1,-2,0,0,1,0,1,1,1,-1,0,0,1,0,0,0,-1,0,-1,0,1,0,0,0,1,1,0,1,-1,2,-1,0,0,0,1,0,1,0,1,-1,-1,0,-1,1,1,-1,-1,0,1,1,0,0,0,1,0,-4,1,0,-1,1,0,-1,1,1,0,2,-3,0,0,1,0,-2,0,0,-1,-1,-1,-1,2,-1,0,2,0,1,1,-1,2,2,1,-1,0,0,1,0,1};
			611: counter1_out = '{0,2,0,0,0,0,2,0,0,1,0,-2,0,-1,0,-1,1,0,0,-1,-2,1,-2,-1,-1,0,0,0,0,-2,0,-1,0,0,0,0,0,0,-2,0,0,1,0,0,1,0,0,2,0,2,-1,0,2,0,1,0,-2,0,0,-1,0,0,1,1,0,1,1,0,-2,0,1,-1,-2,0,2,0,-1,1,2,0,-1,-1,-1,-2,-1,0,1,-1,0,0,0,1,2,-1,-2,1,1,0,0,0};
			612: counter1_out = '{0,-1,0,1,0,0,0,1,-1,-1,0,-1,1,-1,-1,-3,-2,-3,0,-1,1,1,1,0,0,1,2,-1,0,0,-1,0,-1,1,0,2,0,0,0,-1,-1,-2,0,-1,0,0,-1,1,0,1,-1,1,2,0,1,1,0,1,1,1,1,-2,1,0,0,-1,0,0,-1,0,0,0,-1,-1,0,-1,1,1,-1,0,-3,0,-2,1,0,1,0,0,0,0,1,0,-1,-1,0,1,1,0,-1,-1};
			613: counter1_out = '{0,1,0,1,-1,1,1,0,1,0,2,-1,1,-1,0,-1,0,0,1,-1,-1,-1,0,0,-1,2,-1,0,2,-1,2,0,0,1,1,1,-1,1,-1,-1,-1,1,1,-1,-1,0,0,-1,0,1,-1,1,2,0,-1,0,-1,1,0,1,0,-1,-1,0,0,0,0,-1,0,0,-1,0,1,-2,1,0,-2,0,1,-1,-1,-1,1,2,0,0,0,-2,2,1,-2,0,0,-2,0,-1,-1,1,1,-1};
			614: counter1_out = '{1,2,0,1,0,0,0,-1,-3,1,2,2,1,-1,1,-1,-2,3,1,1,-2,1,2,-1,0,0,0,1,1,-2,0,0,0,0,-1,2,1,-2,-1,-2,1,1,0,0,0,-1,-1,-1,-1,2,0,1,0,-1,-2,2,2,2,0,1,-1,0,0,0,-1,-3,0,2,0,2,-1,0,-1,1,0,-1,0,-1,1,-1,-1,2,-1,2,0,0,0,0,0,-2,-1,0,1,0,0,1,0,-1,0,-1};
			615: counter1_out = '{-2,-2,-1,0,1,1,1,0,1,1,1,1,1,-1,0,0,1,2,2,0,0,1,-3,-1,-1,1,-1,0,2,-2,1,1,-1,1,-1,1,0,0,-1,1,1,0,1,-1,-2,0,1,-1,0,0,2,-1,0,-1,0,2,0,-1,1,-1,-1,-1,0,0,0,-2,-2,1,0,0,2,0,-1,1,0,-1,1,-1,1,1,1,0,0,0,-1,1,1,1,-1,1,-2,-2,1,-1,-1,1,1,1,0,-1};
			616: counter1_out = '{-2,-1,1,1,-1,1,1,0,1,-1,-1,0,0,-2,0,0,-1,1,-2,0,2,0,1,0,1,0,-1,1,-1,1,-1,0,0,2,0,0,1,-1,0,1,-2,-1,-1,0,0,-1,-1,0,-2,1,0,-1,1,-1,0,-2,1,-1,1,0,1,1,0,-2,-1,-1,1,0,-1,0,0,0,0,0,-1,1,0,1,0,1,1,1,0,2,0,-1,0,0,0,1,1,0,1,-1,1,-1,0,0,1,-1};
			617: counter1_out = '{0,-1,-1,2,1,-2,0,0,0,1,-1,2,1,-1,0,0,1,0,0,0,1,-1,0,-1,-1,-1,-2,0,1,0,0,0,0,1,-1,0,-2,0,-1,0,0,0,1,0,1,1,0,-1,0,-1,-1,1,-2,0,-1,-2,0,0,0,0,1,1,-1,-1,2,0,1,0,-1,1,0,2,-1,0,-1,-2,-1,1,1,0,0,-1,1,0,-1,1,1,-2,0,-1,0,0,0,1,-2,0,0,-2,-1,-1};
			618: counter1_out = '{-1,0,0,-1,0,0,-1,1,1,0,0,0,-2,0,2,0,1,2,2,0,-1,1,1,-1,0,0,1,1,-1,-1,1,1,0,-1,1,0,-1,1,-1,1,0,1,1,1,2,0,0,-1,0,0,3,-1,0,-1,1,-1,0,1,0,-1,-1,0,-1,-2,0,0,2,0,-1,-1,1,-1,-2,0,1,0,1,-1,0,0,0,0,0,0,1,0,-1,0,1,0,-1,1,-2,0,0,1,1,-1,-2,0};
			619: counter1_out = '{0,1,0,0,0,-1,2,-1,0,1,1,0,-1,-1,2,0,-2,1,-2,0,1,-2,1,-1,1,0,1,-1,0,1,-1,0,-2,-1,0,-1,0,0,1,0,-1,1,1,2,0,-1,1,-1,0,0,-2,0,1,2,-2,1,-1,0,1,0,2,0,-1,1,1,1,0,-1,-1,-1,0,1,0,0,1,-1,1,2,-1,1,0,1,1,0,2,2,0,0,2,0,0,0,1,0,1,-2,-2,0,1,-1};
			620: counter1_out = '{-1,-2,1,-1,0,1,-1,-2,0,-1,0,0,1,-1,0,0,1,-1,0,0,0,-2,2,0,1,0,2,1,1,1,-1,0,-1,0,-1,-1,1,0,-1,-1,0,0,0,0,2,-1,0,0,0,1,1,0,0,0,0,0,0,0,-1,0,-1,0,0,-1,2,-1,0,0,1,2,0,0,1,-2,-2,0,0,1,1,1,-1,0,-1,0,-1,1,-1,0,0,-1,-2,0,-1,0,0,0,0,0,-1,1};
			621: counter1_out = '{2,1,-1,1,-1,-1,0,-1,0,1,0,0,-1,0,0,1,0,1,0,2,1,-1,3,-1,0,-2,-1,-1,1,-1,2,1,1,-2,1,0,0,-1,0,-1,0,-2,1,2,2,-1,2,0,-2,0,-1,1,0,0,-1,-1,-1,0,-2,0,0,-1,1,1,-1,-1,0,0,1,0,0,0,0,1,0,-1,-1,1,0,0,-1,-1,0,-1,-1,-1,1,-1,-1,1,-2,-1,-1,0,0,2,0,0,0,-1};
			622: counter1_out = '{1,1,1,1,0,1,1,1,1,0,0,-1,-1,1,0,0,-2,0,0,0,-1,-1,0,0,0,0,2,0,0,2,1,1,0,2,-2,-1,1,-1,2,-1,0,-1,0,0,-1,0,1,0,2,0,1,-1,1,1,-1,-1,-1,-1,-1,0,0,0,1,2,-1,0,0,2,0,1,-1,-1,1,-1,-1,0,0,-1,-1,-1,-1,0,1,1,-2,-2,-2,0,0,0,0,-1,1,-1,-1,1,1,0,-2,1};
			623: counter1_out = '{0,1,-2,1,-1,0,-1,1,1,0,1,1,1,0,0,2,1,-1,-2,-1,0,-1,1,-1,0,-1,0,0,-2,1,0,3,0,2,-3,0,-1,-1,-1,2,-2,1,-1,-1,1,-1,1,1,0,0,1,-1,0,0,0,-4,1,0,-2,0,-2,-1,-1,1,0,-1,-1,-1,0,-2,0,-1,0,0,0,1,-1,0,0,0,-1,1,1,1,-2,-1,-1,-2,0,0,0,2,0,2,0,-1,0,0,-1,1};
			624: counter1_out = '{2,-1,0,0,1,-2,0,0,0,0,-1,0,1,0,-1,0,-1,0,1,0,0,0,1,-2,1,0,1,0,1,0,1,0,-1,1,-1,0,1,0,1,0,-2,0,1,-1,0,-1,1,1,-1,0,0,-2,0,0,0,1,0,1,-1,1,-1,-2,-1,-2,1,0,0,0,1,-2,-1,-1,-2,-1,1,0,-2,1,0,0,0,0,0,0,0,0,1,-1,0,2,0,0,-2,-1,1,0,0,2,-1,1};
			625: counter1_out = '{-1,1,-3,0,0,1,-1,0,-1,1,-1,0,-2,1,0,0,1,0,0,0,0,-2,-2,1,-1,1,0,0,2,2,0,-1,-1,1,2,0,0,1,3,2,0,0,-1,0,0,1,1,0,0,2,1,0,1,-1,0,-3,-1,-2,0,0,-1,-1,-1,0,1,1,1,0,0,0,0,0,-2,-1,1,-1,-1,1,1,0,0,1,2,-1,1,0,0,-2,0,1,0,1,0,1,-1,0,-1,3,-2,0};
			626: counter1_out = '{0,2,-1,-1,-1,-1,0,1,0,1,0,1,1,-1,0,-1,1,-2,0,0,1,0,0,-2,0,-1,0,0,-1,1,0,0,0,0,0,0,-1,-1,1,0,0,0,1,0,-1,0,1,0,0,0,-1,-1,3,0,-3,-2,1,-1,0,2,1,0,0,0,-1,0,0,0,0,2,1,0,-2,-1,0,-1,0,1,0,0,0,0,1,-1,-1,0,0,1,1,-1,-1,2,-1,0,-1,0,0,0,0,1};
			627: counter1_out = '{1,1,-1,-1,-2,-1,2,1,-2,0,2,1,0,0,2,-1,1,1,1,-1,1,-3,-1,0,2,-1,-1,-1,1,1,1,1,0,-2,1,1,0,0,-1,0,-2,1,1,-1,-3,0,0,0,0,-1,0,1,1,-1,-4,0,1,0,0,-1,-1,0,-1,1,1,1,-1,-1,-1,1,0,-2,1,-1,1,0,1,0,0,2,0,0,0,-1,1,1,-1,-1,0,0,0,0,1,1,-2,1,0,0,0,0};
			628: counter1_out = '{-1,0,1,2,1,0,0,0,2,0,1,1,-1,1,0,0,1,-1,-1,0,0,-1,-1,-2,-1,1,0,-1,1,-1,0,0,1,2,1,0,-1,0,-1,-1,0,-1,-1,0,1,0,-1,-2,0,2,-2,1,1,-1,-2,-2,0,-1,1,0,0,0,2,0,2,1,-1,-2,2,1,0,-1,-1,-1,-1,0,-2,0,-2,0,0,-1,2,0,0,0,2,0,0,1,1,-1,0,1,-2,1,-1,0,1,0};
			629: counter1_out = '{0,1,0,0,0,0,1,1,-1,-2,2,1,-2,0,1,1,2,0,2,0,1,-1,-1,-1,0,0,1,-1,2,0,0,1,-1,0,-1,1,-1,1,-1,-2,-1,2,2,0,-1,-1,-1,1,0,0,-1,1,-1,0,-1,-1,0,0,-1,-1,0,0,-1,1,0,0,1,0,0,1,2,1,-1,1,-1,0,1,2,1,1,-1,0,-1,1,0,-1,0,-1,1,1,1,0,0,1,-1,-2,1,1,0,-1};
			630: counter1_out = '{-1,0,1,2,-1,2,1,0,1,0,-1,1,1,0,0,0,0,1,0,0,-1,-1,-1,1,-1,0,0,-1,-1,-1,-2,0,0,2,0,0,0,1,-1,-1,1,0,0,-1,-1,1,0,-3,1,0,0,1,0,-1,-2,-1,0,1,-1,-2,-2,1,-1,1,-2,1,1,0,0,1,0,-1,1,-1,1,-1,0,1,-1,-1,1,0,0,-2,-1,-2,1,-1,-1,0,0,1,0,-2,-2,0,0,1,0,2};
			631: counter1_out = '{-1,-3,0,0,1,0,0,1,1,0,0,1,-1,1,1,0,0,0,-1,1,-2,0,0,-1,0,0,0,-1,-1,-1,1,-2,0,0,-2,0,-1,1,-1,0,-1,1,0,-1,2,0,0,0,-1,0,0,-1,0,0,-1,0,1,0,0,0,0,0,-1,0,-2,0,0,-1,2,0,-1,0,-1,1,0,0,0,1,0,0,0,-2,0,-2,1,0,0,-1,-1,-2,1,-1,-1,1,0,0,0,0,-1,0};
			632: counter1_out = '{1,-2,0,0,2,0,-2,1,1,-1,-1,0,2,0,0,-1,-1,0,-2,0,-2,2,1,0,1,2,1,1,0,-1,-1,-2,0,1,0,0,-2,1,0,0,0,0,1,0,1,-1,0,1,1,-1,-1,-1,-1,-1,-3,-1,1,0,0,0,0,-1,-1,-1,-2,0,1,1,1,1,-1,-1,0,-1,0,0,-1,0,1,-1,0,-2,0,-1,2,1,2,-1,1,0,0,1,1,1,0,0,-1,1,1,1};
			633: counter1_out = '{0,-1,-1,-2,1,0,0,1,0,-1,-1,-1,1,-1,-1,-1,-1,0,-1,-2,-1,1,0,0,2,0,0,0,0,0,1,-2,-1,1,0,-1,-1,0,0,1,-1,0,2,1,1,0,1,0,-1,1,0,0,0,-1,0,0,-1,0,0,-1,-1,0,0,0,0,1,1,0,1,-1,-1,-2,2,1,-1,2,2,0,1,0,2,-1,-1,1,0,0,0,1,0,0,1,0,1,0,0,0,0,-2,1,0};
			634: counter1_out = '{-1,-2,-1,-1,-1,-1,-1,0,0,-1,-1,3,1,0,1,1,0,1,0,-2,0,0,2,0,-1,-1,0,3,0,0,0,0,0,1,0,0,1,1,-2,-2,0,-1,-1,0,-1,2,-1,1,0,1,-1,-2,0,1,1,0,0,-1,-1,0,-1,-1,0,0,0,0,1,0,-1,-2,0,-1,1,-1,-2,-1,1,0,-1,-2,1,-1,1,-1,-1,0,0,1,2,-3,1,0,-1,0,2,-1,-1,0,-2,0};
			635: counter1_out = '{0,0,-1,-1,-1,-1,-1,2,-1,-2,0,0,0,0,-2,0,0,3,0,0,-1,1,1,1,0,1,-2,0,-1,1,4,-1,1,-1,0,1,1,-1,-1,0,1,3,-2,2,0,-1,0,0,0,1,0,0,-1,1,0,-3,1,0,0,-1,-2,1,0,0,2,1,0,-1,-1,3,0,-1,2,1,0,-1,0,0,0,-1,0,0,-1,1,-3,0,-1,0,0,-2,0,-1,1,0,1,0,1,0,1,-1};
			636: counter1_out = '{1,0,-1,-1,0,0,0,0,-1,1,0,1,1,1,-1,0,0,1,-2,-1,-1,-1,0,0,-1,0,-1,1,0,1,2,0,-1,0,-1,0,-1,1,2,-1,-1,-1,0,-1,1,-1,0,1,-1,1,-2,-2,-1,-1,-1,-1,1,0,1,-1,-1,0,2,-1,1,1,0,0,-1,1,0,0,1,-1,1,-1,-1,-1,1,0,-1,0,-1,-1,1,1,0,0,-1,1,0,-1,-1,-2,1,0,0,1,2,0};
			637: counter1_out = '{-1,0,0,1,0,-2,-1,0,-1,1,-3,1,0,0,-1,1,0,-1,-1,0,-1,1,0,0,2,1,-1,0,1,0,-1,-1,0,0,0,-1,-2,0,1,-1,1,2,-2,0,2,1,1,-1,2,-1,-1,0,0,-1,2,1,0,-1,1,0,-2,0,-2,2,2,1,0,1,-1,-2,0,-2,1,-2,-1,-2,0,-1,-1,0,-2,-2,-1,0,0,-1,0,-1,-1,0,0,2,0,0,2,1,0,-2,0,-1};
			638: counter1_out = '{-1,-1,-1,1,0,0,0,0,-2,-1,1,1,0,1,1,-2,1,0,-1,0,0,0,-1,0,1,1,0,0,-1,1,-2,-1,0,-1,0,1,0,0,0,1,1,0,1,-1,1,0,-1,0,1,0,-1,0,-1,0,0,0,1,-1,2,0,1,1,1,-1,0,2,2,1,0,2,0,-2,-1,-1,-1,1,0,-1,-1,1,0,-1,0,0,1,1,1,0,-1,1,0,-2,-1,-1,-1,0,-1,1,0,0};
			639: counter1_out = '{-1,1,1,1,-2,0,2,0,0,0,-1,0,0,0,0,0,0,-1,1,0,0,0,0,0,-2,-1,1,0,1,1,1,0,1,2,0,-2,0,-1,-2,-1,-1,1,-1,1,1,1,0,-1,-1,0,-1,1,0,2,-1,1,-2,-1,-1,0,-1,0,0,0,-1,0,0,0,-1,0,-1,1,0,0,1,1,0,-1,0,-1,0,0,-1,-1,1,0,1,0,0,0,2,-2,0,-1,-1,-1,0,-1,0,-1};
			640: counter1_out = '{-1,-1,1,0,1,1,-1,0,-2,-1,2,0,2,1,-3,1,1,0,-1,0,1,1,-1,-1,2,0,1,-1,0,0,2,1,0,1,0,1,0,1,0,1,1,-1,-2,0,0,-2,-1,1,-2,0,-1,1,2,-1,2,1,-2,1,0,-1,1,0,-1,1,0,0,0,-1,0,0,0,0,0,0,0,-1,0,1,0,0,-1,2,0,-1,0,-1,0,2,0,-1,1,0,-1,0,-1,0,2,1,-1,-1};
			641: counter1_out = '{0,-1,0,0,1,-2,-1,-1,-1,-2,0,1,1,2,-1,0,1,1,0,-2,-1,-1,-1,-1,0,-1,-1,0,1,-2,0,0,0,0,2,0,1,0,0,0,-2,1,1,0,0,0,1,2,2,1,1,-2,2,0,0,1,1,0,-1,0,0,-1,0,-1,0,0,0,2,0,0,0,2,-2,0,0,0,-1,0,-1,1,2,1,0,-1,1,-1,0,0,-1,0,1,2,0,-1,1,1,2,0,0,1};
			642: counter1_out = '{0,1,-1,1,0,0,0,1,2,-1,0,0,-1,0,-1,0,2,0,0,1,-1,0,1,3,0,0,0,1,0,1,1,0,2,0,1,0,0,2,-1,1,0,0,0,0,-1,-2,2,0,0,0,1,1,1,-1,-1,1,1,1,-2,1,0,0,1,0,-2,-1,0,-1,0,1,0,1,-1,0,2,2,-1,0,1,0,-1,0,0,-1,0,0,0,1,-3,-1,0,-1,1,-2,0,-1,0,1,0,-1};
			643: counter1_out = '{2,0,2,1,-1,0,-1,-1,-1,0,-1,-1,0,1,0,-1,2,0,0,0,0,2,1,0,0,0,-1,1,-1,0,0,0,0,-1,1,0,0,0,0,0,-1,1,-2,0,0,0,0,-1,-1,1,1,0,-1,2,1,0,-1,0,-2,-2,0,0,2,0,-1,0,-1,0,0,0,0,1,-1,0,2,1,0,2,1,-2,0,-2,-2,-1,0,0,3,0,1,1,0,0,1,-1,0,0,-1,0,1,0};
			644: counter1_out = '{-1,-1,-2,0,1,-1,1,-1,1,-1,0,1,-1,1,0,-1,1,1,-1,1,0,-2,-2,-1,-2,0,1,1,0,-1,3,0,-1,0,0,-2,1,-2,0,0,-1,-1,-1,-1,-1,1,2,2,-1,1,-1,-1,-1,0,0,1,-2,1,0,0,0,3,1,1,-1,0,-1,-2,2,2,0,0,0,0,0,1,0,1,-1,-1,1,2,1,-1,2,1,-1,-1,0,1,0,-1,1,0,0,-1,2,-1,-3,-1};
			645: counter1_out = '{2,0,-1,1,0,1,2,0,1,0,1,-1,0,-1,-1,0,1,-1,-2,-1,0,0,1,-1,-1,-1,0,1,-2,0,1,0,0,0,0,1,-1,0,-1,1,0,1,1,0,0,-1,-1,-1,0,0,0,-1,-1,0,-2,-1,-1,0,-1,-1,-1,0,1,-1,1,1,0,0,-1,-3,-1,-1,-1,2,0,0,1,-1,0,-1,1,-1,0,0,3,0,-1,1,-1,2,0,1,0,0,-1,-2,0,1,0,-2};
			646: counter1_out = '{0,1,-2,0,-1,0,-1,1,1,1,0,0,0,0,0,2,0,1,0,-1,0,0,0,0,1,0,0,0,0,0,0,0,1,1,2,-1,1,1,-1,1,0,1,1,1,-1,-2,2,-1,0,-1,2,0,0,-2,-1,1,0,1,2,1,-1,-1,1,-1,-1,-2,2,-2,-1,2,-1,0,-1,1,1,2,0,1,0,-1,0,1,0,-1,0,0,0,0,-1,2,-1,-1,0,0,1,0,2,0,-1,-1};
			647: counter1_out = '{0,-1,-2,-2,-1,-1,0,1,-2,1,-1,-2,0,1,0,-1,0,0,-1,1,0,-1,-1,0,-1,1,-1,-1,-2,0,1,-1,-1,4,1,1,0,0,0,1,0,2,0,-2,0,-1,1,-2,-1,-1,1,2,0,1,0,0,-1,1,1,1,0,0,0,1,-2,1,-4,-1,1,-1,1,1,-2,0,-1,1,-1,0,2,1,1,-1,-1,0,0,0,-1,0,2,0,0,0,0,0,0,-1,-1,1,1,0};
			648: counter1_out = '{-1,1,1,2,0,-2,0,1,0,-2,1,1,2,-1,0,2,0,-1,0,0,0,0,0,-1,1,0,0,0,0,-1,0,1,-2,0,0,-1,0,2,0,0,0,1,0,0,1,0,0,0,2,0,-1,0,0,1,-1,1,1,0,0,1,-2,0,-1,1,0,0,0,0,1,2,1,-1,0,1,0,0,1,0,1,0,0,-1,0,1,0,0,0,1,-1,-1,-1,0,0,0,-1,0,-1,1,1,-1};
			649: counter1_out = '{0,0,0,2,-1,1,0,0,0,-2,0,0,0,0,0,0,1,0,2,-1,0,2,1,0,1,-1,0,-1,1,0,1,0,0,1,1,-1,0,-2,-2,0,0,-1,-1,-1,0,0,2,1,0,-1,-1,0,-1,1,0,0,1,0,0,1,-1,0,0,0,0,0,0,0,0,1,0,-1,-2,1,0,1,1,-1,1,0,0,-1,1,2,-1,1,0,0,-1,1,1,-1,0,0,0,0,1,0,-1,0};
			650: counter1_out = '{-3,1,-2,0,2,0,0,-2,0,1,1,1,1,1,0,1,-1,2,-2,0,1,-1,0,1,-1,0,2,0,1,3,1,-1,0,1,1,-2,1,0,1,0,-1,-1,-1,1,0,1,2,1,0,-1,0,1,0,0,-1,1,-1,2,0,0,0,1,0,0,-1,1,0,1,-1,1,0,0,0,0,0,3,-1,1,1,-2,-1,1,0,-1,-1,-1,1,2,-1,-1,0,-1,1,-1,0,-1,2,-2,-1,0};
			651: counter1_out = '{0,1,-1,0,1,0,0,1,1,1,0,0,0,-1,0,-1,0,-1,-2,1,1,0,0,0,0,0,1,1,1,1,-1,0,-1,-2,0,2,1,0,0,0,-3,1,-2,-3,-1,-2,-2,-1,0,1,0,1,0,2,-1,-1,-1,-1,-1,0,2,-1,-1,-1,1,2,0,2,-1,-1,-1,-1,1,0,0,1,0,0,0,-1,0,-1,3,0,0,1,0,1,-2,1,1,0,-1,-1,-1,1,1,2,0,0};
			652: counter1_out = '{0,0,-1,0,0,1,0,1,-1,-1,3,0,-3,-2,0,-1,0,0,0,1,1,1,-1,0,-1,-1,-1,0,2,1,-1,0,-2,-1,-1,1,-1,0,1,-1,0,0,1,-2,2,0,0,2,-1,0,0,0,1,0,-2,0,0,1,0,0,0,1,0,0,-1,1,0,1,-1,1,-1,-1,-1,-1,-1,0,0,1,1,3,3,1,0,0,0,-1,0,0,0,-2,-1,1,1,-1,0,-1,-1,0,0,-2};
			653: counter1_out = '{-1,0,0,2,0,2,-1,1,-1,2,3,0,0,0,1,0,0,-1,0,0,0,0,1,-2,1,1,0,0,0,0,0,0,0,1,0,1,-2,0,-1,-1,-1,0,0,-1,2,-2,1,0,2,1,-3,-1,-1,1,0,1,0,-1,2,0,-2,1,-1,1,0,0,-1,0,-1,0,-1,0,0,0,2,0,0,0,1,-1,-1,1,1,0,0,0,1,1,1,0,0,0,-1,0,-1,-1,-1,1,1,0};
			654: counter1_out = '{-1,-1,-2,-1,-1,0,1,0,1,-1,1,2,0,0,0,1,1,-1,-1,0,1,-2,-1,0,0,-1,1,0,0,0,1,0,-2,1,0,3,-1,2,2,-1,1,2,-1,0,-2,0,0,-2,2,1,1,0,-1,0,-2,-3,-1,0,3,-2,-2,0,0,0,1,1,0,-3,0,0,1,0,1,0,1,0,0,0,1,1,1,1,1,-1,0,2,-1,0,1,2,1,0,0,1,-1,-1,1,1,0,0};
			655: counter1_out = '{1,0,-1,0,0,0,0,0,0,0,1,0,0,-2,0,0,0,-2,1,0,0,-1,1,-3,0,1,-1,-2,1,-1,2,0,1,0,1,1,2,0,0,0,2,1,-2,0,0,-2,-2,0,-1,1,0,1,2,2,-2,-2,-1,-2,0,0,-3,-1,0,1,-1,-2,-2,0,-1,3,0,2,-1,1,0,1,1,3,0,0,2,0,2,1,1,-1,0,1,0,0,3,-3,2,-1,1,0,1,0,0,-1};
			656: counter1_out = '{0,-1,-1,1,2,1,1,0,1,1,1,1,1,-1,0,-1,-1,-1,1,0,2,0,-1,-1,-2,-1,-1,0,-1,1,0,1,-1,1,0,1,-1,1,0,-1,0,1,0,-2,1,1,1,1,1,0,1,1,-1,0,-2,-1,0,-2,0,1,-1,-1,-1,-1,1,2,1,0,0,0,0,1,0,-1,1,-2,-1,2,2,1,-1,2,1,2,1,-2,-2,0,1,0,2,0,1,1,0,2,-1,0,-1,0};
			657: counter1_out = '{-1,-1,1,0,1,0,2,0,1,0,0,1,1,0,2,-1,0,0,0,0,0,-1,0,-2,1,0,1,-1,-1,0,0,1,0,0,-1,-1,-1,-2,0,2,0,1,-2,0,-1,-1,-2,1,-1,0,-1,0,-1,-3,-2,0,1,-1,1,0,0,1,0,0,1,1,-1,0,0,1,-2,3,-1,2,0,0,0,0,0,1,1,1,3,-1,-1,-1,2,1,0,-1,1,-1,-1,-2,0,1,0,0,0,1};
			658: counter1_out = '{0,0,0,0,0,-1,2,-1,2,0,2,1,0,-2,0,-1,-2,-1,2,-1,0,-1,1,0,1,1,-2,0,1,-1,-1,0,-3,1,0,0,-3,0,0,-2,1,-1,0,2,0,-1,-1,1,1,1,-2,1,1,-1,-1,-1,0,-1,0,1,-3,0,0,0,0,2,0,-2,1,0,1,2,-1,0,0,-1,2,0,1,-1,0,0,1,0,1,-2,0,0,-1,2,3,-1,0,-1,0,0,-1,1,0,0};
			659: counter1_out = '{0,0,0,-1,1,-1,-1,1,1,-1,1,1,-1,-2,2,0,1,1,1,0,-1,0,-1,-1,-1,0,0,0,-1,-1,0,-3,-3,0,0,0,-1,1,-1,0,0,1,0,0,-1,1,0,-1,0,0,1,1,-1,0,1,-1,2,3,-1,-1,-1,0,-1,1,-1,3,0,0,0,-1,1,0,0,-1,0,-1,0,0,2,-1,1,0,2,-2,0,-2,0,0,0,1,2,0,-2,1,1,1,-1,1,1,0};
			660: counter1_out = '{-2,-1,1,-2,-1,-1,2,-1,0,-3,0,0,1,0,2,0,0,1,1,1,-4,-1,0,1,-2,2,0,0,-1,-1,0,-2,1,-1,0,0,-1,0,0,0,0,-1,-2,1,-2,1,-2,-1,1,0,0,0,0,-3,1,0,1,1,-1,0,-2,0,-1,1,0,1,0,1,-1,0,-1,1,0,1,0,3,0,0,0,0,1,-1,2,-1,-1,1,1,0,-1,-1,2,0,1,0,0,0,0,-1,1,-1};
			661: counter1_out = '{0,-2,0,-1,1,-2,-1,0,0,1,0,0,-1,0,1,0,1,2,0,-2,0,-1,-2,1,2,-1,0,-2,-2,-1,-1,0,-1,1,-1,1,-1,1,1,1,0,0,-3,-1,-2,0,1,0,-2,0,-1,0,0,-2,-1,-1,1,-1,0,0,-2,2,0,-1,-1,1,2,1,0,0,-1,0,1,-2,0,0,0,-2,-1,1,1,-1,1,0,1,1,0,0,-1,1,0,0,0,-1,-2,0,0,2,0,2};
			662: counter1_out = '{0,-1,1,0,1,-1,0,0,-1,-1,0,0,0,-2,-1,1,0,-3,0,0,0,0,1,0,1,1,-1,1,1,0,0,0,0,1,1,1,-1,-1,0,2,-1,1,-1,0,0,0,1,2,-1,0,0,1,0,0,0,2,1,-1,-1,0,0,1,0,1,1,2,1,-1,0,0,2,-1,-1,-2,-1,-1,-1,0,1,1,2,2,-1,-1,-1,-1,0,1,0,1,0,0,-1,-1,1,0,0,0,-3,0};
			663: counter1_out = '{0,0,-1,2,-2,-3,1,1,2,-1,0,0,0,-2,-1,0,0,0,-1,-1,0,2,-1,-2,0,1,-1,0,0,-2,0,0,0,0,0,0,1,1,0,2,0,2,0,1,0,-2,0,-2,-1,0,0,0,0,-1,-1,-1,2,1,-2,0,1,-1,-1,0,0,-1,1,2,1,-1,-1,1,1,1,0,2,-1,-2,-1,0,1,0,-2,-2,-1,-1,1,1,2,0,1,0,-1,-1,0,-1,-1,1,-1,0};
			664: counter1_out = '{-1,1,0,-1,-1,0,-1,0,0,0,0,2,-1,0,-1,0,-1,-1,0,-2,-1,2,-1,0,-1,0,0,0,-2,-1,0,-2,0,0,-1,-1,1,0,0,0,-2,1,-1,2,1,-2,1,1,-1,0,-2,1,0,-1,-1,-2,-2,0,1,-3,1,-1,2,-1,-1,1,0,0,-1,0,1,-1,1,-2,1,1,0,0,0,0,1,3,0,0,0,2,0,0,0,1,1,-1,-1,0,0,1,0,0,-2,1};
			665: counter1_out = '{0,1,0,1,-2,-1,-1,2,1,-1,2,-1,0,-1,-1,0,0,1,0,-1,-1,0,1,1,-2,1,-1,1,-1,-2,-2,0,0,1,1,-1,1,-1,-1,0,1,0,-1,0,1,1,0,-1,-1,0,1,1,-1,-2,-1,-1,0,-1,0,0,-1,0,2,-1,2,1,-1,0,1,-1,1,1,-1,-4,-2,0,-1,0,-1,1,0,-1,-1,-1,-2,0,-1,0,0,0,2,0,0,1,0,2,1,1,0,0};
			666: counter1_out = '{2,1,1,0,-1,0,1,0,0,1,0,-1,1,0,2,0,0,-1,-1,0,0,0,1,-1,0,1,0,-1,1,0,1,2,2,-1,0,-2,1,-2,1,0,-3,1,-1,0,-1,0,1,1,0,0,-2,-1,0,-2,2,1,1,0,1,1,1,-1,-1,0,0,1,0,-1,-1,-1,-2,1,0,2,-2,-1,1,1,0,1,-1,0,0,2,0,0,0,1,-1,-1,-2,0,-1,1,-1,1,-1,1,0,-2};
			667: counter1_out = '{-1,1,2,0,0,-1,2,1,-1,3,-1,1,-1,0,-1,0,0,1,1,0,0,0,1,-3,-1,0,1,0,-1,0,0,2,-2,-1,1,1,0,0,0,1,2,1,0,0,1,1,-1,0,0,1,-1,0,-1,3,1,0,0,0,0,1,-1,1,0,0,-2,0,0,0,-2,0,1,-1,0,0,0,0,-1,0,0,-1,0,2,-1,1,0,1,0,3,1,-1,-1,-1,1,0,-1,1,-1,0,0,2};
			668: counter1_out = '{0,1,0,0,0,0,1,-1,1,0,2,0,-1,-1,0,0,0,1,0,-1,1,0,2,-1,0,-1,0,-1,0,-1,0,0,-1,2,-1,0,0,-1,-2,-2,0,1,-1,-1,-1,0,0,0,0,0,0,1,1,1,2,0,-1,-2,1,-1,2,-1,0,1,1,0,1,0,0,-1,2,0,2,0,1,1,2,0,1,1,1,1,0,2,1,1,1,0,1,-2,0,0,2,-1,1,0,1,1,-1,0};
			669: counter1_out = '{-2,0,0,-1,0,-1,-2,0,-1,-2,1,1,-3,-1,0,1,-1,1,1,-1,-1,0,-1,0,1,-1,1,0,1,0,0,0,0,-3,0,-1,-3,1,2,0,1,0,0,0,0,1,1,1,-1,-1,-1,0,0,0,0,-3,0,-1,-1,1,-2,-1,1,-2,-1,0,-1,1,-1,-2,1,1,0,-1,0,-1,0,0,1,0,0,0,-1,1,0,0,1,0,0,-1,0,1,0,0,-1,0,0,0,0,-1};
			670: counter1_out = '{1,0,2,-1,2,-1,0,2,1,0,0,-1,-1,1,0,-4,1,-1,-1,1,0,-1,-1,2,0,-1,0,0,-2,0,-1,1,-1,1,-1,1,0,1,0,0,1,1,0,1,-1,0,-1,-1,0,-1,0,0,0,0,1,0,-1,1,-1,0,-1,-2,0,1,-2,0,0,1,1,-2,-1,-1,0,-1,0,0,0,2,0,0,2,0,-1,0,0,0,-1,-2,-1,0,0,1,0,-1,-2,-1,-1,0,-1,0};
			671: counter1_out = '{1,0,1,0,0,0,0,-2,-1,0,-2,-2,0,-1,0,-1,0,-2,1,1,0,1,1,-1,1,0,2,0,0,0,0,0,1,-1,-1,1,-1,1,0,0,-1,2,-1,0,-2,0,1,0,-1,0,-1,0,1,1,0,0,3,-2,-1,1,1,-1,-2,1,-1,2,0,-1,1,1,1,0,2,1,2,1,-1,-1,-1,0,0,0,1,0,1,-1,1,-1,0,0,2,-2,2,-1,-1,2,0,1,-1,-1};
			672: counter1_out = '{1,0,0,0,0,-1,1,2,-1,2,0,-1,-1,1,-1,0,1,1,0,0,0,0,-1,1,0,0,0,0,0,-1,0,0,-1,0,0,0,2,0,1,0,1,-1,1,-2,-1,-1,0,-1,1,-1,-1,0,0,-2,0,2,0,0,2,0,0,1,0,0,0,0,-1,1,0,0,1,-1,0,0,0,-1,2,0,-1,-1,0,-3,-1,0,-2,-1,-2,1,0,-1,1,1,0,1,1,-2,1,1,0,2};
			673: counter1_out = '{1,0,0,2,-1,0,-1,0,-1,-1,0,-1,-1,0,-1,1,1,-1,1,-1,-1,-1,0,-1,-1,1,0,-2,1,-1,0,-1,-1,-1,-1,1,3,0,1,1,0,0,-2,0,1,1,1,0,-2,0,0,0,0,1,-2,1,-2,-1,1,-2,0,0,0,-1,-1,1,-1,0,0,0,0,1,-1,1,-1,0,0,0,0,0,0,-1,0,2,-2,1,0,-1,0,-2,0,0,-1,1,0,0,0,1,0,1};
			674: counter1_out = '{1,1,0,-1,0,-1,0,0,0,-1,0,0,-1,1,0,1,1,2,0,0,0,-3,0,1,1,0,1,-1,-2,0,1,0,0,-1,0,-1,0,-2,1,0,2,1,0,-1,0,-2,0,-1,0,1,1,1,2,0,2,1,2,0,1,1,0,-1,0,1,0,1,0,1,0,0,0,0,-2,1,1,0,-1,-1,2,0,0,0,0,-1,-1,0,0,2,0,0,0,-1,1,0,-1,0,-1,-2,0,0};
			675: counter1_out = '{-1,0,1,1,0,1,0,0,-2,-1,0,1,1,-1,1,2,0,-3,-1,1,1,0,1,0,4,1,2,-2,0,0,-1,1,0,2,1,-1,1,1,1,0,3,2,1,0,-1,1,0,-1,1,0,0,0,-1,0,0,0,0,0,0,0,1,-1,0,1,-1,-2,1,-2,-2,0,1,-1,0,-1,0,1,0,1,1,1,0,0,1,-1,1,1,-1,0,3,-1,1,-2,1,-2,-1,-1,1,0,1,-3};
			676: counter1_out = '{1,0,0,0,1,0,0,0,0,-1,-1,-1,1,1,-1,-1,-1,0,-1,2,1,0,1,0,0,-1,0,1,1,-1,-1,1,1,0,0,1,2,0,-1,0,0,0,0,0,0,-1,-2,0,0,0,0,1,0,0,-1,0,-2,0,1,0,0,0,0,-1,1,-1,0,0,0,-1,0,-1,1,-1,0,0,0,1,-1,-1,0,1,-1,0,1,-2,-1,1,-1,1,0,1,0,-2,0,0,0,1,1,0};
			677: counter1_out = '{0,3,1,2,-1,1,-1,-2,-1,-1,-1,-2,1,1,0,-2,-3,0,-1,0,1,0,0,2,1,0,-3,0,3,0,1,0,-3,1,1,0,2,-1,0,2,2,2,-1,0,-1,0,-1,1,-1,0,0,-2,1,1,0,-1,2,-1,0,1,1,0,1,-1,2,1,-1,1,0,-1,0,-2,0,0,-1,-1,0,0,1,1,-2,-2,0,0,-2,0,0,-1,-1,0,0,2,-1,0,2,-1,-3,0,1,0};
			678: counter1_out = '{0,0,0,0,0,3,0,0,0,0,2,-1,0,-1,1,1,0,1,-1,1,1,-1,0,0,3,0,-1,1,-1,2,2,1,-2,0,1,1,0,3,1,-2,0,-2,-2,-2,0,1,0,-1,0,1,1,0,0,-1,-2,-1,0,-1,0,-1,1,0,0,-2,-1,-1,0,0,-2,-2,0,0,1,0,0,0,1,-1,1,0,1,1,-1,-2,-3,1,1,-1,2,0,-1,1,1,0,0,0,1,0,2,1};
			679: counter1_out = '{-1,0,0,0,1,3,0,1,0,2,-1,1,0,0,2,0,-4,2,-1,-1,1,-1,1,0,2,-1,-2,2,2,0,0,1,0,-1,2,0,-1,-1,0,-1,-1,0,-1,1,-1,1,-1,1,1,0,2,1,-1,0,0,-1,1,1,-1,0,1,-3,2,1,0,0,-1,1,-1,2,0,-1,-1,0,2,0,1,2,2,-1,0,1,-1,-1,-1,0,0,0,-1,0,0,1,-1,1,-1,1,1,0,0,0};
			680: counter1_out = '{-2,0,0,-1,0,-1,0,0,0,2,-1,1,0,1,0,2,-1,-1,-2,0,0,0,1,0,0,1,1,-1,1,1,2,-1,0,1,-1,0,1,1,-1,-1,-1,1,0,-2,-2,3,-2,1,1,0,1,-1,0,-1,-2,1,0,0,0,0,0,-1,1,-1,-2,-2,1,1,-2,1,-1,-1,0,0,-1,0,0,-1,0,0,1,0,1,-2,0,-1,1,0,1,0,0,1,-1,-1,0,-1,-3,-1,1,0};
			681: counter1_out = '{0,1,-1,-1,1,-1,-1,0,0,1,1,1,1,-1,0,0,-2,0,-1,1,1,-2,0,0,-1,-1,1,0,0,0,2,2,1,0,-1,2,1,0,0,0,0,-3,0,-1,0,-1,-1,0,1,1,-1,-1,-1,-1,-3,0,2,1,-1,-1,1,-1,1,-1,-1,1,0,0,1,1,0,1,-2,-2,0,0,1,0,1,-1,0,0,-1,1,-1,0,0,-1,1,-2,1,0,0,-1,0,1,1,0,0,0};
			682: counter1_out = '{-1,-2,0,1,-1,-2,-1,-1,0,-1,1,-2,0,0,2,1,1,1,0,-1,-2,2,0,0,1,0,1,0,1,0,1,0,0,-1,-1,2,0,-1,0,0,1,-1,0,-1,-1,2,0,0,-2,-2,0,1,0,1,-1,-2,1,-1,0,0,-1,-1,0,0,-1,0,0,0,-1,0,1,-1,-2,-1,2,1,0,0,0,1,1,1,-1,0,-1,2,1,0,2,-1,2,0,0,-1,1,1,0,-1,2,0};
			683: counter1_out = '{-1,1,0,0,1,1,1,0,1,1,1,0,0,-1,1,-1,-1,1,0,1,2,-1,-1,-2,1,-1,0,2,0,1,-1,0,0,-2,1,0,0,0,1,1,1,0,-1,-2,0,1,0,-2,0,2,0,1,1,-2,-1,0,0,0,0,2,0,1,0,-1,-1,-1,1,-2,0,-1,1,0,0,-1,0,0,0,0,0,-3,0,0,-1,-1,2,1,2,-1,1,0,1,-1,0,-1,0,1,1,0,-1,1};
			684: counter1_out = '{1,-2,-1,1,0,1,0,-1,0,-1,0,1,1,-1,0,0,0,2,1,0,1,0,-1,0,0,0,0,0,0,0,1,-1,-1,0,-1,0,0,1,0,-1,-1,-1,-2,-1,0,-1,0,2,0,-1,-1,-1,1,0,-1,0,0,0,-1,1,1,-1,-1,0,-1,-1,2,0,1,-1,1,0,1,-1,-1,0,1,-1,1,0,1,-2,0,0,0,-3,-2,-1,1,-1,1,1,-2,0,0,1,0,-1,1,0};
			685: counter1_out = '{-1,-1,-1,1,-1,0,0,0,2,0,2,0,-1,0,0,0,1,2,-1,2,0,0,-1,0,0,0,0,1,0,1,-1,2,1,1,1,2,0,1,0,-1,0,-1,-2,0,-1,-1,-2,-1,1,1,0,1,0,0,-3,0,-1,-2,0,0,-2,-2,-2,-1,-1,-1,0,-1,0,0,-1,0,-3,0,0,1,0,2,0,-1,0,0,0,-1,1,-1,1,-1,0,0,1,-1,0,0,0,-1,0,-1,1,1};
			686: counter1_out = '{1,-1,-1,1,2,1,1,1,2,0,3,2,-1,-2,1,1,-1,-1,0,1,-1,2,0,-2,1,0,0,0,-1,-1,-1,1,-1,-2,1,2,0,0,0,-2,0,1,-3,0,-3,-1,1,0,-1,2,0,1,0,0,0,0,0,2,1,-1,-3,2,0,1,-1,0,0,-1,0,0,1,0,0,0,0,0,0,0,0,0,1,1,0,0,-1,0,1,0,-1,1,0,0,-1,-1,-1,2,-1,0,0,0};
			687: counter1_out = '{0,0,-1,-1,0,0,1,0,0,-2,0,1,0,-1,1,-1,1,1,0,1,-1,-1,1,0,-2,1,1,0,0,-2,0,1,0,0,0,1,-1,0,0,0,1,1,-1,-2,0,3,-1,-1,0,0,0,-1,-1,0,-4,-1,1,0,1,1,-2,0,-1,0,1,-2,0,-1,2,1,0,-1,1,2,0,-1,-1,1,-1,0,0,0,1,-1,1,0,0,0,0,1,-1,-1,1,0,-1,0,-1,1,0,0};
			688: counter1_out = '{-1,-1,0,1,0,1,-1,-1,0,-1,-1,1,1,1,2,-1,-1,2,-2,0,-1,1,-1,0,0,-1,-1,1,-1,-2,1,-1,-1,1,1,-1,-1,0,1,-1,-1,2,1,1,2,-1,0,-2,-1,1,1,-1,-1,-1,1,0,1,1,-1,-1,1,-1,0,0,0,0,0,-1,-1,0,1,2,1,-1,0,0,0,0,-1,-1,0,1,-1,-1,1,-1,-1,1,1,-1,1,1,2,-2,1,2,1,1,0,-1};
			689: counter1_out = '{-1,0,2,-1,0,-1,-1,2,1,1,2,0,-1,0,1,0,1,0,-2,-1,-3,0,-1,0,3,1,1,0,0,0,-1,1,1,1,1,1,-1,0,0,1,1,1,-1,0,0,2,-1,2,0,1,-1,1,-1,0,3,-1,1,1,-1,0,-1,0,-1,1,-1,1,0,0,-1,-1,0,-1,0,0,-2,0,2,-1,2,-1,1,1,-1,-1,-1,-1,0,1,0,1,0,-1,-1,0,0,0,2,0,0,-1};
			690: counter1_out = '{-1,2,-2,1,0,-2,1,1,0,0,1,1,-2,0,0,-1,-1,-1,1,0,-1,-2,-1,-1,-1,-1,-1,-1,0,-3,-1,1,-1,-1,-1,0,-1,-1,1,2,0,0,-1,-2,1,1,0,0,1,0,0,-1,-1,-1,1,-2,-1,0,0,1,-1,-1,-1,3,1,1,1,1,2,-2,1,-1,-1,0,1,0,1,-1,-2,0,2,0,-1,0,1,2,0,-1,-1,0,1,-1,1,-2,-1,0,0,0,0,0};
			691: counter1_out = '{-1,0,3,0,-2,-1,0,0,-1,2,0,1,-1,0,1,0,0,0,-1,1,0,2,0,0,0,-1,0,0,0,0,0,-1,2,-1,1,-1,0,0,2,1,-2,1,0,1,1,0,2,-1,0,-1,0,-1,-1,1,-2,-1,2,0,2,0,-1,1,0,0,2,1,0,-1,1,-3,1,0,-1,0,0,1,3,0,-1,1,3,0,-1,-1,-2,1,-1,1,0,1,0,1,2,-1,0,-1,0,0,0,1};
			692: counter1_out = '{1,-2,1,0,0,0,1,-1,0,2,0,0,1,-1,0,0,0,0,-2,-1,0,0,0,1,0,0,1,1,0,0,-1,0,1,0,0,0,1,-1,1,0,-1,1,-2,-1,1,2,-1,-2,0,0,-1,1,0,-1,1,-1,0,-1,1,0,0,0,-1,-1,1,0,1,0,0,0,0,0,0,-1,0,0,1,0,-1,-1,0,0,-1,-1,0,1,-1,0,-3,1,-1,-1,1,-1,1,-1,-1,-2,1,0};
			693: counter1_out = '{2,1,1,0,-1,0,1,1,0,1,0,-2,2,-1,0,-2,0,1,0,0,-1,-1,1,0,1,1,0,0,1,0,0,1,0,-1,-1,-1,0,0,0,0,0,-1,-1,-1,0,1,0,1,0,-1,-1,0,0,-1,0,1,0,1,0,-1,0,-2,1,-1,1,-1,-1,-1,-1,-1,0,-1,0,-1,0,0,0,-1,0,-2,2,1,1,0,1,1,0,1,0,-1,-1,-1,0,-1,0,1,1,0,0,-1};
			694: counter1_out = '{-1,0,2,0,-1,0,0,-1,1,0,0,0,1,-1,0,0,0,0,0,0,-1,-1,1,-3,-2,0,0,1,1,0,-1,1,-1,0,0,1,0,-1,-1,1,-1,-2,0,-1,-1,0,2,0,-1,0,-1,0,-2,2,1,0,-1,0,0,0,0,0,0,0,0,-1,2,-1,2,0,0,0,0,1,1,1,1,1,1,-3,1,1,-2,1,0,0,-3,0,0,1,1,-2,-1,1,1,1,1,0,2,1};
			695: counter1_out = '{-1,0,-1,0,1,-1,2,0,-1,1,0,-1,2,0,-1,0,0,1,1,0,1,0,0,-1,1,-1,-1,0,1,0,1,0,2,-2,-3,-1,1,0,-1,0,2,0,-1,1,0,1,-1,0,1,0,0,0,-1,-2,1,-1,0,2,-1,-1,-1,0,-2,-2,-1,1,-2,-1,1,1,2,0,-1,1,-1,-2,2,0,-1,0,0,0,1,-1,0,0,0,0,-1,0,-1,-1,0,1,-2,2,0,1,-2,0};
			696: counter1_out = '{-2,0,-1,-1,0,0,1,2,0,0,-1,-1,0,0,0,1,0,1,0,0,1,-1,0,2,2,0,-1,-2,0,-1,-1,0,1,0,1,0,1,0,-1,0,-1,-2,-1,1,1,-1,2,0,-2,0,0,0,-1,0,0,-1,0,0,-1,-1,1,0,-2,-1,0,1,0,1,0,1,0,1,0,1,1,0,-1,1,1,0,-1,0,0,0,-1,1,1,0,1,-1,1,1,2,-1,0,-1,-2,0,-1,-2};
			697: counter1_out = '{0,2,0,0,-1,1,0,-1,-2,-1,-1,-2,1,0,0,-2,0,-1,1,-1,0,-2,1,0,-1,-1,-1,2,0,1,0,0,-1,0,2,1,2,2,-1,0,0,-1,0,-1,0,1,2,-1,0,2,-1,-1,-1,1,1,0,0,-1,1,-1,0,-1,-2,-1,0,-1,0,-1,-1,1,0,0,2,0,2,1,1,0,0,-2,0,-1,-1,0,1,1,1,-1,1,0,0,1,-1,0,0,1,0,0,2,0};
			698: counter1_out = '{1,0,0,-1,-1,0,0,1,0,1,-1,1,-1,-1,2,0,0,-1,1,0,0,0,-2,-1,0,2,0,0,1,0,0,0,0,0,-1,-2,-2,2,0,-1,-2,-1,0,0,0,0,0,1,-1,1,1,-1,1,2,0,1,0,0,1,0,-1,3,0,0,0,-1,0,1,-3,-1,0,0,-1,0,1,0,0,1,-1,0,-1,0,-2,0,0,2,0,0,0,0,2,-1,1,0,0,-1,0,1,1,-1};
			699: counter1_out = '{-1,2,1,0,1,0,-3,0,0,-1,1,0,0,1,-1,0,0,0,0,-1,1,-1,3,-1,0,-1,0,1,-1,1,0,1,1,-1,1,1,-1,-1,1,2,1,0,-1,0,0,0,0,0,1,1,-1,0,-1,-1,1,0,0,0,0,1,-2,-1,0,1,0,0,-1,0,2,0,1,1,2,1,0,0,0,0,-3,0,0,0,0,1,-1,0,-1,1,0,1,1,0,0,0,-1,1,0,1,1,0};
			700: counter1_out = '{-1,1,1,-1,-1,-1,-1,1,1,1,0,-1,1,-1,2,-1,0,-1,1,1,1,-1,-1,1,-1,0,0,-2,0,2,-1,-1,0,0,1,1,-1,2,0,0,0,-1,1,0,1,-1,1,1,-1,1,1,0,0,0,-1,2,-1,1,0,-2,1,1,1,-1,2,0,2,0,-2,1,-2,0,0,1,0,0,-1,1,0,1,1,0,0,0,0,-2,0,1,1,2,0,1,0,1,-2,-1,2,-1,0,0};
			701: counter1_out = '{2,0,0,-1,1,1,-1,0,-1,-1,-1,-1,-2,1,1,0,0,-1,-2,0,1,-1,0,-1,0,-1,0,0,0,1,0,1,1,2,0,0,0,0,-1,1,-1,-1,1,2,1,0,1,0,0,1,-1,0,1,0,1,-1,0,1,-1,0,0,1,-1,0,0,-1,1,-1,1,1,0,0,-1,0,0,-1,-1,-1,0,0,1,-1,-2,0,0,-1,0,-1,0,-2,0,-1,-1,0,0,-2,0,0,1,0};
			702: counter1_out = '{-1,0,1,0,0,0,0,-1,-2,1,-2,0,1,1,1,0,1,0,0,-1,0,0,0,0,1,1,-1,-1,1,1,1,-1,1,-1,-1,1,-1,1,1,1,0,0,-1,0,0,-1,0,-2,1,1,-2,-1,1,1,1,1,0,0,0,0,0,0,1,-1,0,1,-1,-1,0,-1,1,0,-1,-2,0,-1,1,1,-2,0,-1,0,0,-1,0,-2,-1,1,2,-1,1,0,-1,1,0,-1,1,1,0,1};
			703: counter1_out = '{0,0,-2,-1,0,-3,2,-1,0,-2,0,1,0,0,1,-1,0,-1,0,-1,0,0,0,-1,-2,1,1,-2,0,-1,0,-1,-1,0,-2,-1,0,2,1,1,1,-1,1,2,-1,2,1,0,0,-1,-1,0,0,0,-1,0,0,0,0,0,-1,0,1,2,0,1,-1,1,-1,1,1,0,-2,1,-2,-1,0,-2,-1,0,1,0,1,-1,-1,1,2,0,0,0,-1,-2,2,-1,0,-2,-1,-1,-2,0};
			704: counter1_out = '{0,1,2,-1,-2,-1,2,1,-1,1,0,1,0,-1,0,0,0,-1,1,1,0,1,0,0,-1,1,-1,0,1,1,0,2,1,0,1,1,0,2,0,0,-1,0,1,-3,-2,0,0,0,0,-1,0,0,-1,1,-1,0,0,0,2,-1,0,-1,-1,-1,1,0,-1,0,1,0,0,-1,1,0,0,1,1,0,0,1,0,-1,-1,1,-2,1,1,-1,0,2,-2,-1,0,1,-1,-1,0,-2,2,-2};
			705: counter1_out = '{0,1,1,0,0,-1,1,1,-1,1,0,1,-2,0,0,-1,-1,0,0,2,1,1,-1,0,1,0,-1,-1,0,1,1,0,1,-1,-1,-1,2,1,2,0,1,1,0,-1,0,1,-1,-1,0,-1,-2,1,-1,-1,2,0,0,1,0,1,0,-1,0,-1,0,-1,0,1,0,0,0,-1,-1,1,-1,1,0,-1,-2,1,-1,0,-2,0,0,1,1,1,1,0,0,2,1,-1,-2,-2,1,1,2,1};
			706: counter1_out = '{1,-1,1,0,0,1,-1,0,0,-1,0,0,1,0,1,1,-1,-1,0,0,0,1,-2,0,2,1,1,1,0,-1,1,1,0,1,0,-1,-1,1,1,-1,-2,-1,0,0,1,1,-1,0,0,0,2,0,-1,2,0,0,2,-2,-1,-1,-1,-1,1,-1,0,-1,1,-1,0,1,0,1,0,-1,-1,-2,0,1,1,2,1,0,-1,1,-2,0,-2,1,-1,-1,0,0,0,1,0,2,1,-1,2,1};
			707: counter1_out = '{2,-1,2,0,0,1,2,-1,-1,-1,0,1,0,0,1,0,-1,-2,-1,-2,1,-2,0,-1,0,0,1,-1,2,0,1,1,-1,-1,-1,-2,-1,1,0,1,0,2,0,-1,0,2,0,-1,1,0,0,0,0,1,-1,0,-1,2,-1,-1,1,-2,0,0,-1,1,1,1,0,1,-2,-1,-2,-1,0,-1,-1,-2,0,0,0,0,-1,0,-1,1,1,-2,-1,-1,0,0,-1,1,0,-1,2,-2,0,1};
			708: counter1_out = '{0,0,0,-2,0,1,1,1,0,-1,0,1,-1,2,0,0,-1,0,0,0,0,2,0,-1,0,-1,0,-2,0,0,1,-1,-1,0,1,1,2,1,0,-1,0,1,1,0,0,0,1,1,1,0,1,0,-2,0,0,0,2,1,2,0,-2,-3,0,-1,0,0,-3,-1,1,0,0,0,0,0,-1,0,-1,1,1,-1,-2,-1,0,0,1,-1,1,1,1,0,0,-1,-2,0,1,-1,-1,0,-1,-2};
			709: counter1_out = '{0,0,1,2,-1,-1,0,2,0,-2,1,-1,0,-4,0,1,1,1,0,-2,0,0,0,-1,1,-1,-2,2,-2,-1,0,-3,0,-2,1,1,1,1,1,-1,3,-1,-1,-1,0,0,1,-1,0,-2,1,0,-1,-1,-1,-1,0,2,-4,0,2,0,1,0,-2,-1,2,1,-1,-1,1,1,1,-1,-2,0,1,1,-1,-1,-1,0,1,-1,-2,2,0,2,2,0,1,-1,-1,-2,-1,0,2,0,1,1};
			710: counter1_out = '{0,-1,-1,1,0,3,0,0,3,0,0,-1,1,1,0,1,2,0,-1,0,-2,1,2,-2,1,-2,-2,0,0,-2,2,3,0,0,0,0,-1,1,0,0,1,1,0,-2,0,3,-1,1,1,1,1,1,-1,0,0,-1,-2,0,0,-1,0,1,-1,0,0,-1,1,0,-1,1,0,-1,-2,1,-2,1,1,1,-1,-1,-2,-1,0,-1,0,0,0,2,1,-1,-1,1,-1,-1,0,1,-1,1,-1,-1};
			711: counter1_out = '{1,1,2,1,-1,-1,-1,0,3,-1,0,0,1,2,1,2,2,1,0,0,-1,1,0,-1,0,1,1,0,1,0,0,1,-2,0,1,0,1,-1,0,-1,1,0,-2,0,1,0,-1,-1,-1,0,3,0,-1,-1,1,-1,0,0,-1,0,1,1,-1,0,0,-1,1,0,0,-2,-1,2,1,1,-1,1,-1,1,1,0,0,1,1,-3,1,1,0,0,0,-2,-1,0,0,-2,0,2,1,-1,0,-1};
			712: counter1_out = '{-2,0,0,1,0,2,0,-3,2,0,1,1,1,1,1,0,1,-2,-1,0,1,2,0,-1,-1,0,0,0,1,-2,-1,-1,0,3,1,2,0,-1,-1,-2,0,-1,0,0,1,0,0,0,1,-1,3,0,1,1,0,-1,1,2,0,2,0,-2,-1,0,0,-1,1,1,0,0,0,2,0,1,0,-1,-1,1,1,2,-2,0,0,0,3,0,1,0,-2,1,1,-1,-3,-2,1,1,1,0,-1,-1};
			713: counter1_out = '{1,0,1,1,-2,0,-1,-1,1,0,-1,2,-1,0,0,1,0,1,0,0,0,0,0,0,0,0,-2,-1,0,-1,-1,2,1,-1,0,0,0,1,1,0,2,-1,-1,-2,0,2,-1,0,0,1,0,-1,-1,-1,1,1,0,0,1,1,-2,0,0,-1,-2,0,-1,0,0,1,-1,1,2,-1,0,0,1,-2,0,1,-1,-1,0,1,0,-1,0,0,-1,0,0,0,1,0,1,-2,0,1,0,0};
			714: counter1_out = '{-1,-1,0,0,-1,-1,0,-1,1,0,1,0,-1,1,-1,1,0,1,0,1,0,1,-1,0,-1,1,0,-1,0,-1,-2,1,-1,1,-1,0,-2,1,1,2,2,-2,-1,1,1,1,0,1,1,2,3,-1,0,1,0,-1,1,2,1,0,0,-1,0,0,-1,-1,-1,0,0,-1,0,-1,1,1,-2,0,0,0,0,-1,-2,-1,0,0,-1,0,-1,0,-1,-1,2,0,0,-1,-1,1,0,-1,-1,0};
			715: counter1_out = '{-2,0,2,0,1,0,0,-1,0,-1,0,0,-1,0,-1,0,2,0,2,-1,-2,1,0,0,-1,-2,1,0,-1,-1,1,-1,-1,1,-1,0,1,2,-1,-1,2,-1,-1,0,0,0,0,-2,1,0,1,1,1,-1,1,1,2,0,1,0,0,1,-1,-1,2,0,0,0,1,0,0,-1,0,1,0,0,0,-1,0,2,0,-1,-1,0,0,0,-1,0,-1,1,1,0,-1,0,-1,1,0,-1,-1,1};
			716: counter1_out = '{-1,0,-1,1,0,-2,1,0,1,1,-1,0,0,-1,0,0,0,-1,1,2,-2,2,0,-2,0,1,-1,0,2,2,1,0,-1,-1,-1,1,-1,0,1,2,-1,-1,-3,0,-1,0,0,1,2,-1,1,0,1,-1,0,0,1,3,0,1,1,-1,2,-1,0,1,0,1,0,1,-1,-1,-2,1,0,0,1,0,-1,-1,0,1,0,0,-1,1,0,0,-1,0,0,1,-1,-1,0,1,0,0,1,1};
			717: counter1_out = '{-1,2,1,1,-1,-1,1,-1,0,1,-1,2,1,0,1,1,-1,1,1,1,-2,0,0,-2,0,1,0,0,-1,-1,1,-1,-1,0,0,0,-1,0,0,0,0,-1,-2,-2,-2,1,1,-1,1,0,2,0,-1,1,1,-1,1,3,0,-2,0,0,-1,1,2,2,1,1,1,-1,-1,0,0,2,-3,0,0,-1,0,0,1,1,0,1,0,2,0,1,0,-1,-2,-1,1,-1,-1,1,0,1,1,0};
			718: counter1_out = '{-1,-1,1,-1,1,-1,-1,0,2,1,1,0,0,0,1,0,0,-1,0,0,0,2,-2,-1,-2,1,2,2,0,0,0,-1,0,-1,1,0,1,1,-1,1,-1,-1,-1,-2,-1,1,1,1,0,-1,2,-1,0,-1,1,-2,-2,2,2,-2,1,-1,1,-1,1,2,2,0,-1,1,-2,0,0,0,-1,-1,1,-1,0,-1,1,1,1,0,0,1,0,1,1,2,-1,-1,1,-1,1,-1,1,1,0,1};
			719: counter1_out = '{-1,1,0,-1,1,-1,2,0,0,-1,1,-1,0,1,1,-3,-1,0,0,-1,0,1,-1,0,0,0,0,-3,-3,0,0,0,0,0,0,-2,-2,-1,2,0,-1,1,0,-2,1,0,1,-1,-1,0,-1,1,-2,0,-2,-2,1,0,-1,0,1,1,0,-1,1,1,0,-2,1,0,0,1,1,0,0,0,1,0,1,-2,1,0,-1,0,0,-1,-1,2,-1,-1,-1,0,1,-1,0,1,0,-1,1,0};
			720: counter1_out = '{0,0,1,-1,0,-2,1,0,0,0,-1,0,0,1,-1,-1,2,-1,0,-1,0,0,0,2,0,1,0,-1,0,0,-1,1,1,0,-1,-1,1,-1,1,0,1,-1,0,-2,0,1,0,-1,-1,0,1,0,0,0,1,-2,1,0,1,0,-1,-1,0,-1,0,2,-1,0,-1,0,-1,-1,-2,-1,-1,0,1,1,1,-1,2,1,-1,0,1,1,-1,0,-1,2,2,0,1,-2,1,1,0,-1,0,0};
			721: counter1_out = '{0,0,0,-1,1,1,2,0,2,0,0,0,1,-2,1,1,1,0,0,-2,0,0,-2,0,0,-1,-1,-1,1,0,1,1,0,-1,1,2,0,1,1,1,-1,0,1,1,1,2,0,0,-1,0,2,2,0,0,1,0,0,1,-1,0,-1,1,0,0,1,0,1,3,-1,1,3,0,-1,0,0,-2,0,0,-1,0,0,1,-1,0,2,1,0,1,0,1,1,0,0,-1,0,-1,0,-2,-1,0};
			722: counter1_out = '{0,1,1,0,1,-2,-2,0,-1,0,-2,0,0,-1,1,0,-1,1,1,-1,0,1,0,1,-2,0,0,1,1,-1,2,-1,2,1,1,0,0,0,1,-1,0,-1,0,0,1,-2,0,0,2,2,-1,-2,0,0,0,-1,0,0,1,0,0,0,-1,0,-1,2,-1,0,-1,-3,0,0,2,-3,0,0,0,0,-1,0,0,1,0,1,0,0,0,-1,-1,2,1,0,0,0,1,0,-1,1,0,0};
			723: counter1_out = '{3,-3,-1,-1,1,0,0,0,1,0,-1,0,-1,0,0,-1,0,1,0,0,-1,1,0,-1,0,-2,0,0,-1,-1,-2,2,2,-2,0,2,1,0,1,1,1,-1,0,0,0,0,0,-1,0,-2,0,0,-1,0,0,-2,0,1,0,-1,0,-1,0,0,-2,0,-1,0,0,-2,0,0,0,-1,-1,1,0,0,1,1,0,-1,-2,-2,1,0,0,0,0,0,0,-1,-1,0,0,0,0,-1,-1,-1};
			724: counter1_out = '{0,0,0,1,-1,1,0,0,0,1,0,1,0,0,0,0,-2,0,1,1,0,0,-3,0,0,-1,2,-1,-1,-1,-3,1,0,1,-1,-1,-1,0,1,-1,0,2,0,-1,1,-1,0,0,-1,0,1,0,0,0,-1,3,1,1,0,1,0,0,0,-2,0,0,0,1,-2,-1,1,0,1,-1,0,0,0,0,0,-2,0,1,-1,0,0,-1,-1,0,0,0,-1,-2,0,0,-1,2,-1,0,1,0};
			725: counter1_out = '{-1,1,-1,-1,1,-2,1,0,2,1,0,0,-2,1,0,-1,-1,1,1,0,-2,2,-1,0,1,1,0,-1,-1,0,0,1,-1,-2,-2,-1,0,1,-1,1,0,-1,2,-1,-1,1,-2,0,0,-1,1,0,-2,0,0,1,-1,-2,-1,1,-1,0,0,-1,1,0,-1,-1,1,0,1,0,0,-1,2,-1,0,1,-1,0,-2,-1,0,2,-1,0,-2,-2,-1,1,0,-1,1,1,1,-1,-1,-1,-1,-1};
			726: counter1_out = '{0,0,1,0,1,0,1,0,0,0,0,-1,-1,-1,0,2,0,0,1,0,0,0,1,1,-2,0,1,0,0,0,1,0,0,1,-2,0,-1,0,0,-2,1,1,0,-1,1,1,2,0,-1,1,1,0,0,-2,0,-1,1,2,0,0,-1,1,0,-1,0,0,0,-1,2,-2,0,-1,-1,1,-1,0,0,1,1,-1,0,1,0,1,-1,1,-2,-1,1,-1,0,-2,-2,0,0,1,0,0,1,0};
			727: counter1_out = '{1,0,1,0,2,2,0,2,1,0,0,1,0,-2,0,1,0,0,-1,0,0,0,0,-2,-2,0,3,1,1,1,-1,3,-1,0,-1,-1,0,0,2,0,1,-1,0,3,-1,0,0,0,-2,-1,-1,-1,0,1,1,0,-1,1,-2,0,0,-1,1,-1,0,0,1,1,-2,-2,-1,0,-2,-1,0,0,-1,0,0,-1,0,0,0,0,0,1,2,0,0,0,1,0,1,0,-1,-2,2,0,0,0};
			728: counter1_out = '{1,0,1,-1,1,1,0,0,0,0,1,-1,2,1,-1,0,0,-1,0,2,0,0,1,-2,-1,-1,0,-1,3,-1,-1,0,0,-1,0,0,1,0,-1,0,-1,-1,1,2,2,0,0,0,2,1,-1,0,0,2,1,1,1,-3,2,0,0,1,0,-1,-2,0,1,0,0,-1,-1,0,-1,1,-1,1,1,-1,0,-1,0,0,2,-1,0,0,3,-2,-1,-1,0,0,1,-1,-2,-1,1,1,-1,-3};
			729: counter1_out = '{1,-2,0,2,1,1,1,-1,-1,1,0,1,1,0,0,2,0,-2,1,1,1,-1,1,-1,-1,1,0,-1,1,0,-1,-1,0,1,-1,1,1,1,0,0,-1,0,1,1,0,0,1,-1,-1,0,1,-1,0,1,0,1,0,1,1,0,-1,0,1,-1,0,0,-1,1,-2,-1,1,0,-2,1,0,0,1,0,0,1,0,1,2,-1,1,-1,1,1,-1,0,1,0,-2,0,1,-1,0,-1,1,0};
			730: counter1_out = '{-1,1,1,0,0,0,-1,-1,-2,0,0,-1,-1,-1,1,0,0,0,-1,0,1,1,-1,-2,-2,0,-1,1,0,-1,-1,-2,-1,1,-1,2,1,0,0,0,0,2,0,1,1,1,1,-1,0,-1,-1,-1,1,1,0,0,0,0,1,-2,1,-1,0,0,1,1,1,-1,0,-1,1,-1,0,-1,2,1,1,0,2,-1,1,1,-1,-1,1,-2,0,-1,0,-1,-2,0,-1,2,0,-2,1,0,0,0};
			731: counter1_out = '{-1,0,-1,2,0,0,1,-1,0,0,0,-3,-1,-1,1,1,-1,0,-1,0,0,0,-1,1,-3,0,-1,-3,0,1,-1,-1,-1,0,1,0,-1,-1,1,0,1,-1,1,0,0,0,-1,-1,-1,2,-1,1,-1,0,0,1,-1,-1,-1,1,-1,2,-1,-2,-1,-1,0,0,-2,-1,0,1,-3,-2,0,0,1,1,0,-1,2,-1,1,-1,-1,0,2,0,0,-1,0,-2,-1,0,-1,1,0,0,-1,0};
			732: counter1_out = '{-1,0,0,0,0,-1,1,1,-1,1,0,1,-2,0,-1,0,-1,0,2,-2,1,0,-1,-1,0,1,1,1,0,0,-1,-2,0,-2,1,0,-1,1,2,1,0,0,-1,0,-1,0,0,0,1,0,-2,-1,2,0,-2,0,1,-1,1,0,1,0,-1,-2,-2,0,2,-1,0,1,-1,-1,-1,0,-1,0,0,0,-1,2,0,1,0,0,-1,0,1,0,0,-1,-1,1,-1,0,2,0,-1,2,1,0};
			733: counter1_out = '{1,1,-1,0,1,0,-1,1,-1,0,0,-1,-1,-2,-2,0,-1,-1,1,0,-1,0,-1,-1,0,0,-1,1,1,0,2,0,1,-1,-1,-1,1,-1,-1,1,2,0,1,1,-2,0,1,-3,1,0,0,1,0,-1,0,1,1,0,1,2,0,1,0,-1,-1,-2,1,-1,-1,0,-1,-1,0,0,1,1,1,0,-1,0,-2,0,2,-1,0,-1,0,-1,1,0,2,-1,0,0,1,1,0,1,0,3};
			734: counter1_out = '{0,-1,1,0,0,0,1,1,0,1,-1,0,0,-1,0,-1,-1,0,1,0,1,-1,0,-1,0,0,-1,0,0,2,0,-1,2,-1,-1,-1,-1,0,0,-3,-2,0,-3,1,-1,0,0,-1,1,1,0,0,-1,1,-1,1,-2,-1,0,0,0,1,-1,1,-1,-1,0,0,-1,0,1,-1,2,-1,2,-1,0,-2,0,2,0,1,1,-1,1,1,-3,2,-2,1,0,-2,-1,-1,0,-1,-1,0,0,-1};
			735: counter1_out = '{-2,0,-1,0,1,-2,0,-1,-1,1,-1,2,0,1,-2,1,0,-1,1,-1,-1,-3,0,3,-1,-1,-1,0,2,0,0,0,-1,-2,0,-1,0,0,0,2,1,0,-1,1,0,-1,1,0,-1,-2,1,0,0,0,1,0,0,-2,-1,-1,0,-1,-2,0,0,-2,0,0,-1,1,1,-1,1,-1,0,-1,-1,-1,-1,0,1,0,-1,-2,-2,1,-2,1,0,1,-1,1,-1,-2,-1,0,-1,0,1,1};
			736: counter1_out = '{0,-2,0,0,-2,1,0,0,-1,2,1,1,1,0,0,-1,-1,1,0,1,0,-1,-1,0,-1,1,-1,0,-2,-2,0,-1,-1,1,1,0,0,-1,0,1,-1,-1,0,1,1,0,2,-1,1,0,0,-1,-2,-1,-1,1,1,1,1,0,1,1,-2,0,-1,-1,0,0,1,0,1,0,0,1,0,0,0,1,0,1,-1,0,0,0,1,-1,-1,1,1,0,0,-1,-1,1,-1,-1,1,1,1,1};
			737: counter1_out = '{1,0,1,0,0,-2,-1,1,0,1,-1,1,0,0,0,-1,0,1,0,-2,1,0,-1,1,0,1,1,1,1,1,0,1,0,1,-2,0,0,-1,-1,0,2,-1,-1,-2,1,0,1,-2,0,-1,2,1,1,3,-2,-1,-1,1,-1,0,1,0,1,1,0,-1,1,0,-1,0,0,-1,1,2,0,1,0,0,0,0,0,3,1,-1,0,-1,2,0,0,-1,1,0,0,-1,1,0,-1,-1,0,1};
			738: counter1_out = '{1,-2,0,-1,0,0,0,1,1,1,-1,0,1,0,-1,0,-1,-1,0,0,0,2,-1,-1,-1,1,0,-1,-1,2,2,-2,-1,1,-1,3,0,-2,-1,-1,-2,-1,-1,-1,0,0,0,-1,0,-1,1,2,1,1,0,-1,0,1,0,0,1,1,1,0,1,1,1,-1,1,1,0,1,0,-1,0,1,0,-2,0,-2,0,0,-1,0,-1,2,0,-1,0,1,-2,0,0,-2,-2,1,1,0,-1,1};
			739: counter1_out = '{0,1,0,0,-1,1,0,0,0,0,-1,1,-2,-1,2,-2,-2,1,2,1,-1,0,0,0,1,0,0,-1,-1,0,1,0,3,-2,1,-1,1,-1,-1,0,0,0,0,0,-1,1,0,0,0,1,0,-1,0,-1,2,0,-2,0,0,0,1,-1,-1,0,-1,0,-1,-1,0,-1,1,0,0,-1,1,0,2,-2,2,0,0,0,0,2,-1,0,-1,0,-1,1,1,0,0,-2,0,1,0,1,1,0};
			740: counter1_out = '{-1,-1,1,2,0,1,0,1,-1,0,-1,2,-1,-1,0,-1,0,-1,1,1,-1,0,-1,1,-1,-1,1,0,0,1,-1,1,1,0,-1,0,-1,0,-1,0,-1,-1,-1,-1,1,2,-1,-2,-1,1,-1,-2,0,-1,1,-3,0,0,0,0,0,1,0,2,0,-1,1,-2,-2,0,0,0,0,-1,1,0,2,1,-1,0,0,-1,0,-1,0,-1,0,0,0,2,0,-1,0,-1,1,0,0,0,0,0};
			741: counter1_out = '{0,-1,0,-1,0,1,1,1,0,-1,1,2,0,-1,2,0,0,-1,-1,0,0,1,1,1,-2,-1,1,-1,0,2,1,1,1,0,-1,-1,1,0,-1,0,2,0,-1,-2,-1,0,0,-1,0,-2,0,-1,1,0,0,0,1,0,-1,-1,1,1,-1,-1,0,0,0,1,0,0,1,1,-1,0,0,1,0,0,0,0,0,2,-1,0,-1,-1,0,-1,0,2,1,1,1,-1,0,0,0,1,-1,1};
			742: counter1_out = '{1,0,0,0,-1,1,1,-1,0,-1,1,0,-2,0,0,0,0,-3,-1,-2,1,1,1,1,-1,1,0,-2,0,-2,-1,-1,2,1,1,-1,0,0,0,0,1,-2,-1,0,3,1,0,1,0,-1,0,-2,0,0,-1,0,0,-1,0,0,-1,0,0,-1,0,0,2,1,-1,0,3,-1,-1,0,0,-2,1,0,-2,1,0,0,0,-1,0,0,0,-2,1,0,1,2,2,-3,0,1,-3,-1,0,0};
			743: counter1_out = '{-1,0,1,0,-1,1,-1,2,-1,-1,0,0,0,0,0,-1,-1,-1,0,0,0,0,-1,0,1,0,0,0,1,0,-1,1,1,-1,1,0,-1,0,-1,0,-1,-1,1,1,-1,0,1,0,0,1,0,-1,0,1,-1,-1,1,0,-1,-1,1,-1,-2,0,0,-1,-1,1,-1,0,0,1,-1,-2,1,2,0,0,0,1,1,0,2,1,1,1,-1,-1,-1,0,1,0,2,-1,0,1,-1,-1,-1,0};
			744: counter1_out = '{1,1,0,2,0,-1,1,0,0,2,0,1,0,1,-1,0,-1,-1,0,0,0,0,0,-2,0,1,-1,0,-2,1,0,-1,0,0,-1,0,-1,0,-1,3,1,-2,0,0,2,1,1,0,0,0,2,0,0,-1,0,-2,1,0,-2,0,1,-1,-1,-1,1,0,1,0,-2,1,-1,1,2,-1,0,1,0,1,-1,1,-2,0,1,-1,2,-1,1,0,-1,1,0,1,2,-1,2,1,1,1,0,0};
			745: counter1_out = '{0,0,0,0,-2,0,0,1,0,1,-2,-1,1,0,2,1,0,0,0,1,0,2,0,0,1,0,-1,-1,0,-2,-1,-1,0,0,-1,1,-1,0,1,1,-1,-1,-1,1,1,1,0,-1,0,2,1,-2,0,0,-1,0,-1,-1,2,0,-1,-1,1,0,0,0,2,-1,1,2,0,1,-1,1,0,-1,1,0,-1,0,1,3,1,0,-2,0,1,0,1,-1,0,0,0,-1,1,0,-3,-1,0,1};
			746: counter1_out = '{2,1,1,0,0,2,0,1,-2,-1,-1,-2,-2,0,1,-1,0,0,1,1,0,2,1,1,1,0,-1,-1,-1,1,-2,0,1,1,-1,1,-1,-1,0,0,1,-1,0,-2,-1,1,0,-1,2,2,1,0,-1,-1,-1,0,-1,0,0,0,1,-1,2,-1,0,1,0,1,0,1,-2,1,0,1,-1,0,-1,0,2,-2,1,1,1,-3,1,-1,0,-1,-1,-1,0,0,0,0,2,2,-2,-1,-1,1};
			747: counter1_out = '{0,-1,0,-1,0,1,1,1,0,0,0,0,1,-1,-1,1,-2,2,1,0,-1,-1,-1,0,-1,-1,0,1,-1,-1,-1,1,0,0,0,-1,0,0,-2,1,0,1,-1,1,0,0,-1,1,1,0,1,0,-1,0,3,-1,0,0,1,1,0,-1,1,1,0,1,1,0,2,1,0,-1,1,-2,0,-1,-2,0,-1,0,-2,0,1,1,0,-1,1,0,-1,-1,1,-1,0,-1,1,1,0,0,-2,1};
			748: counter1_out = '{-1,0,1,0,1,1,0,3,0,0,0,1,-1,2,0,0,0,-1,-3,1,-1,0,2,-1,-1,0,0,0,-1,-2,-1,0,-1,0,-1,1,0,1,1,0,2,-2,-1,-2,1,0,1,0,-1,1,2,0,0,-1,0,1,1,1,0,-1,0,-1,-1,0,-1,1,1,-1,1,0,1,2,1,0,-1,0,0,0,0,1,1,0,-1,0,0,0,0,2,1,1,-1,-1,-1,0,-1,0,0,0,0,-1};
			749: counter1_out = '{0,0,-2,-1,0,0,-3,-1,-2,0,1,-2,1,0,-1,0,2,0,0,0,1,-1,1,-1,-1,-1,1,-1,1,0,0,0,-1,-1,0,0,-2,0,-1,-1,-1,-1,0,1,1,1,-1,1,1,-3,1,0,-1,1,-1,-1,-1,-1,0,-1,1,-2,-2,-1,1,1,-1,0,0,0,0,0,0,1,1,1,3,-2,-1,0,-1,1,0,0,2,0,0,0,0,1,-1,-1,0,0,-1,-1,-2,1,-1,0};
			750: counter1_out = '{1,0,-2,-1,-1,0,0,1,-2,-1,1,2,-1,-1,1,2,-1,-1,1,0,1,0,0,-2,0,-1,1,0,-1,-2,-2,-1,1,-1,-1,0,-1,0,-1,-1,1,-2,-1,-1,-2,-2,0,0,1,0,0,0,0,0,1,1,0,0,-1,2,1,-1,0,-1,-1,-2,-1,-1,0,0,1,1,0,0,1,0,0,1,1,-1,-1,0,-1,1,0,0,0,-1,0,-1,0,-1,0,1,1,0,1,-1,-1,1};
			751: counter1_out = '{2,1,0,0,-1,0,0,-1,1,2,1,-1,-1,0,1,1,0,0,0,1,0,-1,-1,0,1,1,-1,0,0,0,-1,0,2,-2,1,-1,1,-1,-2,1,2,-1,1,0,1,0,0,0,0,0,2,-1,0,1,0,1,0,1,-1,0,0,-1,1,1,0,-1,0,1,0,1,0,1,-1,0,0,-1,0,-1,1,-2,0,0,-1,-1,0,1,0,1,0,0,0,1,0,-1,0,-1,-1,1,-1,-1};
			752: counter1_out = '{0,1,-1,2,0,1,3,0,1,0,0,-3,-2,1,0,1,0,1,1,0,-1,0,2,0,-1,0,1,1,-1,0,2,0,-1,2,0,-2,-1,0,-1,-1,0,-2,0,-2,1,1,-2,-2,1,-1,-1,0,1,-1,-2,-2,0,0,-2,1,1,0,-1,1,1,1,2,1,1,0,0,1,0,1,0,1,-1,-1,0,0,0,-1,1,-1,1,1,0,0,-1,1,3,0,-1,-1,0,1,-1,0,-2,-1};
			753: counter1_out = '{1,-4,0,1,0,0,0,0,0,1,1,0,0,0,0,0,0,2,0,1,0,0,-2,-1,1,0,0,0,1,0,2,-1,0,0,1,1,1,0,-1,0,0,0,0,0,0,2,-2,0,0,0,-1,-2,1,2,-1,1,1,0,1,1,0,1,0,1,1,-1,-1,0,0,-1,0,0,2,0,0,-2,-1,1,1,0,0,-1,-2,-1,0,0,-1,-1,0,1,1,0,2,0,-1,1,2,3,-2,-1};
			754: counter1_out = '{0,0,1,0,-1,0,0,1,1,0,1,3,1,-1,0,-1,0,1,0,-1,1,0,0,-1,2,-1,0,1,-1,1,0,-1,0,0,-1,-1,0,-3,-1,0,0,0,-1,0,0,-1,1,0,-1,0,1,-1,2,0,-1,0,1,1,-1,-2,-1,-1,1,0,0,0,-1,-1,0,-1,1,-1,-1,1,1,-2,2,1,1,-1,-1,-1,1,-1,1,-1,1,1,1,0,0,1,0,-1,-2,0,0,0,-2,0};
			755: counter1_out = '{0,2,2,-2,0,-1,1,0,-1,0,1,0,0,-1,0,-1,0,-1,0,1,-1,0,-1,0,0,0,0,1,0,1,0,2,1,-1,0,1,1,0,1,1,0,1,0,0,0,1,1,0,2,0,0,0,0,1,-1,-1,-2,-1,-2,-1,2,0,1,0,0,0,-1,1,0,0,0,1,-3,0,-2,0,1,0,1,0,0,0,1,-1,0,0,0,-1,0,1,0,-1,0,1,0,-1,0,-1,0,1};
			756: counter1_out = '{-1,0,-1,-1,1,-1,1,0,0,0,1,1,1,0,0,1,0,0,-1,2,-1,1,1,1,1,2,0,0,1,2,1,0,1,0,1,-2,1,0,1,0,-1,2,0,1,-1,-1,-1,-2,0,1,2,0,1,-2,0,-2,1,0,-1,2,-1,-1,1,-2,-1,1,2,-1,-1,-1,0,1,1,-1,1,2,1,0,-1,1,1,-1,0,-1,-1,-1,-1,0,0,0,0,0,0,0,-3,0,-1,1,1,-2};
			757: counter1_out = '{0,0,-2,0,-1,1,-2,2,-1,1,1,-2,-1,1,1,1,0,0,0,0,-1,-1,0,-2,1,0,2,1,-1,0,-1,0,-1,0,2,-1,1,1,-1,-1,-1,-1,0,0,-1,-2,-1,-1,-2,0,-1,0,-1,0,1,0,1,0,1,0,0,-1,0,-1,0,2,0,0,1,0,-1,-1,2,1,0,0,0,0,0,-1,-1,1,0,0,1,-1,0,1,0,1,-1,0,0,0,-2,-1,0,0,1,0};
			758: counter1_out = '{-1,1,1,0,1,0,-2,1,-1,0,-1,0,0,2,-1,2,2,0,-1,-1,-1,0,1,0,1,0,0,-1,0,0,0,-1,1,0,0,1,0,-1,0,0,1,-2,0,1,-1,0,-1,1,-1,0,0,-2,2,0,0,0,0,1,0,1,1,0,-2,-1,-1,0,1,1,0,1,1,0,-1,-1,1,0,-1,1,0,2,1,-3,-2,0,1,1,0,1,1,0,0,1,0,0,0,0,0,1,-1,0};
			759: counter1_out = '{1,0,1,0,0,0,0,-1,-1,-1,1,0,-1,0,1,0,0,1,3,1,0,-1,0,2,1,-2,-1,-1,-1,-1,-2,-1,-1,1,0,2,-2,0,0,0,-1,0,0,-1,1,0,0,1,-1,0,1,0,0,0,0,-2,1,-1,0,0,0,2,-2,0,0,1,0,1,-2,-1,-1,-1,0,0,-1,0,1,-2,1,1,0,-1,-1,1,0,1,-1,1,0,0,1,0,1,1,1,0,0,0,-1,1};
			760: counter1_out = '{0,0,0,0,0,1,-1,0,0,-2,-1,0,1,1,0,-1,0,-2,-1,0,-1,2,0,0,0,-2,-3,-1,-1,-1,0,1,-2,0,-1,0,0,1,0,-2,-1,0,0,2,1,0,-1,1,-1,0,-1,-1,-1,0,1,1,-1,-1,-2,-2,1,0,1,1,0,1,-1,0,0,0,0,1,0,-1,1,0,1,1,0,1,-1,-1,-1,-1,-1,-1,1,0,0,-1,1,1,-1,-1,-1,-1,0,0,-1,0};
			761: counter1_out = '{0,-1,0,1,1,-1,0,-1,1,0,0,0,0,0,2,1,0,1,1,0,1,0,1,-1,-2,1,-1,1,0,1,1,-1,1,0,1,-1,2,1,-1,1,-1,0,0,1,1,-1,0,-1,0,0,1,0,2,0,1,-2,-1,1,1,-1,2,-1,0,0,1,0,-1,1,0,0,1,-1,1,-1,0,-1,-1,1,0,3,0,0,-2,1,-1,0,-1,1,0,-1,-1,3,0,0,0,1,0,0,0,-1};
			762: counter1_out = '{-1,-1,0,1,-2,-2,1,-2,2,1,0,1,1,-1,1,0,1,-3,0,1,0,0,0,0,2,1,-1,-2,2,-1,1,0,1,0,0,1,1,-1,1,-1,0,2,0,1,0,0,1,-1,0,-2,0,0,-1,-2,1,-1,0,0,-3,0,0,0,-1,-1,-2,2,-1,1,1,0,1,0,-1,0,1,-1,3,1,-2,1,1,0,0,0,1,2,1,0,0,-1,-2,0,-1,1,-3,0,0,-1,1,-1};
			763: counter1_out = '{1,1,-1,1,0,-1,0,1,0,1,1,0,0,-1,0,-1,1,1,3,-1,0,-1,1,0,0,0,0,-1,0,1,0,2,1,-1,0,0,0,1,0,-1,0,0,-1,-3,1,1,0,0,1,-2,-1,1,0,-1,1,-1,1,-1,-1,1,-2,1,2,0,-3,-3,-1,0,-1,0,1,-1,2,0,-1,-1,-1,-1,0,0,-2,-2,-2,1,0,0,2,-1,0,-1,1,-1,-1,0,0,1,0,-1,-1,-1};
			764: counter1_out = '{1,0,2,-1,-1,0,1,0,0,2,-1,2,-2,0,0,1,1,-2,1,0,0,0,1,1,1,1,0,2,0,0,-1,-1,-1,0,1,1,0,-1,1,0,0,-1,-2,0,0,1,0,2,0,-1,1,0,2,0,-1,2,1,0,2,0,0,1,1,2,0,2,0,1,0,0,1,0,0,-1,0,0,1,0,-1,0,-2,-2,1,-2,-2,0,0,-2,2,1,-1,0,-1,-1,0,0,0,0,1,0};
			765: counter1_out = '{1,0,1,-1,0,1,0,0,-1,-1,1,0,1,0,-1,0,-1,0,1,0,-1,0,1,1,1,-1,-1,1,-1,1,0,-1,1,0,0,-1,-1,0,-1,0,0,0,1,2,0,1,-1,-1,0,0,1,0,0,-1,0,3,2,0,0,0,1,0,-1,1,-1,0,-1,-1,2,0,1,1,1,1,1,0,0,0,-2,1,0,0,0,-1,-1,-1,-1,1,1,0,1,0,1,-1,0,0,0,-1,-1,2};
			766: counter1_out = '{0,0,0,0,0,1,0,1,-3,-1,1,1,1,0,0,0,0,0,0,1,-1,-1,0,-1,-1,1,-1,0,-1,-1,0,-1,0,2,1,0,0,-2,-1,0,-1,0,1,1,-1,0,-1,-1,1,0,0,2,0,0,-1,1,0,-1,0,0,0,-1,0,-1,0,0,1,0,-1,0,1,0,0,1,-2,1,0,1,1,0,-2,1,0,-1,1,0,0,-1,0,1,1,-2,-1,0,2,2,-1,-1,1,-1};
			767: counter1_out = '{0,0,0,0,1,2,0,2,0,-1,0,1,0,1,0,2,1,0,0,0,0,0,0,1,1,-1,2,1,2,1,1,1,-1,1,-1,0,-1,0,2,1,-1,0,-1,-1,-1,0,-1,-1,-1,-1,1,0,0,0,1,-1,0,-1,1,-1,-2,1,0,-1,-1,0,2,0,0,0,0,0,-1,0,-1,1,0,2,-1,-2,1,-1,0,0,1,0,0,-2,1,0,0,-1,1,1,1,0,0,-1,1,1};
			768: counter1_out = '{2,0,0,0,1,-2,0,1,0,1,1,3,0,1,-1,0,-1,0,-1,2,0,0,1,-1,1,0,-1,0,-1,0,1,-1,0,-1,0,-2,1,-1,1,-1,0,-2,1,-1,-1,0,3,-1,-1,1,3,0,-1,-1,0,0,0,-1,-1,1,-1,-1,0,2,1,0,0,1,1,0,-1,3,1,0,1,-1,1,0,1,0,-1,1,-2,1,0,-1,-2,-1,-1,1,0,0,1,1,0,0,1,-2,-1,-1};
			769: counter1_out = '{-1,0,1,1,0,0,2,0,0,1,-1,-2,0,1,-1,-1,0,2,0,0,0,0,0,1,0,0,1,-1,0,0,0,2,0,0,0,1,1,0,2,1,-1,-1,0,0,0,0,0,0,1,1,-1,0,0,1,1,0,-1,1,0,0,1,1,2,1,-1,1,-1,0,0,-1,1,1,1,2,0,0,0,1,0,0,2,-1,-1,1,2,0,0,-2,0,1,1,-1,-1,0,1,1,-1,0,0,0};
			770: counter1_out = '{-1,0,0,1,-1,0,-1,-1,-1,0,0,-1,1,0,-2,0,1,-1,1,1,1,-1,-1,0,-1,1,0,-1,-2,0,0,1,-1,-1,-1,3,0,-2,-1,-1,0,0,0,-2,-2,1,0,1,1,0,-1,2,-1,-1,1,0,0,0,-1,0,1,1,0,0,-1,0,-1,-2,0,-2,0,2,0,-1,0,-2,-1,0,-1,-2,0,0,0,-1,-1,-1,0,1,2,0,0,0,0,2,1,0,0,0,1,-2};
			771: counter1_out = '{1,2,0,-1,-2,0,-2,1,0,0,-2,-1,1,1,0,1,0,1,0,0,-1,1,-1,-1,1,-2,0,1,0,-2,0,-1,0,0,0,1,0,-4,0,0,1,0,-2,0,-1,-1,0,-1,-2,2,-1,1,1,0,1,0,-1,0,0,0,1,0,0,-1,-1,2,0,0,1,1,0,1,1,-1,0,-1,-1,0,-1,-1,-1,-1,-1,1,1,0,1,0,1,1,0,-2,2,1,0,0,-1,1,1,1};
			772: counter1_out = '{-1,0,0,0,-1,1,0,0,-1,1,-1,1,1,-1,1,0,-2,1,1,1,0,0,1,0,1,1,2,-1,1,1,1,-1,2,0,-1,0,0,2,-1,-2,-2,-1,-1,0,0,-1,0,0,0,-1,-1,-2,1,0,-1,-1,0,1,0,0,-1,0,-1,1,1,1,0,0,1,2,-1,0,-1,1,-2,0,-2,0,1,0,0,0,1,-1,-1,-1,0,0,0,-2,0,-1,-1,2,0,1,1,-2,-1,-1};
			773: counter1_out = '{1,0,-2,-1,-1,-1,0,-1,1,1,1,0,0,-1,-1,1,2,0,0,0,0,0,2,-1,-1,-1,1,-1,-1,-1,-1,-1,0,0,2,-1,-1,0,1,1,-1,0,1,-2,0,-1,-1,0,-2,1,0,0,-1,-2,0,-2,0,0,0,0,-1,-1,0,0,-2,-1,-1,-3,0,0,0,2,-1,1,-1,2,1,0,-2,0,-2,2,0,-1,1,0,1,0,0,0,0,-2,-1,0,-2,0,-2,-2,2,0};
			774: counter1_out = '{-1,1,2,-2,0,-1,0,0,-1,0,0,0,-2,0,0,-1,3,-1,0,-1,1,0,0,0,1,2,0,0,1,1,-2,-2,1,0,0,0,-1,0,0,-1,2,0,-1,-3,0,0,0,-2,1,-1,0,0,-3,0,1,2,0,0,2,0,0,0,-1,0,1,1,-1,0,1,-2,-2,0,0,0,0,1,0,-1,1,0,1,-2,0,-1,0,-2,2,-2,0,0,-1,-1,0,-1,0,0,2,1,0,2};
			775: counter1_out = '{0,-1,1,1,1,1,1,-1,0,-1,2,1,0,0,1,1,1,-2,0,1,-1,2,-2,0,0,0,2,0,-1,2,1,-1,0,0,-1,-1,-2,-1,-1,1,1,-1,1,-1,0,0,0,-2,2,1,1,-1,1,0,0,-1,1,0,0,0,3,0,0,0,-1,-1,0,0,1,-1,0,1,-1,0,1,-2,1,-1,-1,0,2,1,0,0,-2,0,1,1,0,-1,-2,1,1,0,1,-1,2,-1,0,-2};
			776: counter1_out = '{2,0,0,0,1,-1,-1,0,-2,1,0,0,-1,0,1,-1,0,0,0,1,0,1,-1,1,-3,0,0,-1,1,0,-1,-1,0,-1,-1,-1,2,1,1,1,1,0,1,1,1,1,1,0,0,0,0,1,1,0,0,-1,-2,0,1,1,-1,1,1,-1,1,0,-1,2,0,1,-1,0,0,0,-1,2,0,1,0,0,1,2,0,-1,0,-2,1,0,2,0,2,0,1,0,0,-1,-2,-2,0,0};
			777: counter1_out = '{-1,0,1,1,0,0,1,0,-1,-1,0,-2,-1,0,1,0,0,1,0,0,0,0,0,1,0,1,0,0,0,1,-1,1,-1,2,-1,-1,0,-1,2,-1,0,-2,0,-1,0,-1,1,-1,1,-1,-2,0,0,1,0,1,2,-2,0,0,0,-2,0,-1,1,3,1,0,1,1,0,1,0,-1,0,1,-1,-2,0,0,1,2,-1,0,-2,0,-1,0,0,0,1,1,0,-1,-2,0,0,1,1,0};
			778: counter1_out = '{-1,0,0,0,1,0,0,1,0,3,0,-1,-2,-1,0,1,-2,-2,1,-1,-1,-1,1,1,0,0,0,0,-1,0,-1,1,1,-1,3,1,2,1,-1,0,0,0,1,0,-2,2,0,1,0,0,1,1,1,0,0,1,0,1,0,0,0,0,0,0,1,1,0,0,0,-1,1,0,2,1,0,0,1,-1,2,0,1,-1,0,-1,1,0,0,1,1,2,0,0,0,1,-1,0,0,0,0,0};
			779: counter1_out = '{1,0,0,-1,2,-1,-1,1,-1,0,0,0,1,-1,0,0,1,0,-1,0,0,1,0,1,0,1,-1,-3,-1,0,0,0,-1,2,1,-2,0,1,-2,0,-1,1,-1,0,-1,2,-2,1,1,1,-1,-1,0,-2,0,0,1,0,1,0,-1,0,1,1,0,1,0,0,0,-1,2,0,-1,2,-1,-1,0,0,1,-1,-1,1,-2,-1,-1,1,0,0,0,1,-1,0,0,-1,0,0,0,-1,1,-1};
			780: counter1_out = '{0,2,-1,0,0,0,-3,-2,0,0,-2,1,1,-2,0,0,0,-1,0,0,1,-1,1,1,2,0,-1,1,-2,0,0,0,1,0,-1,-1,0,0,1,-1,1,0,-1,1,-1,2,-2,0,0,0,-1,1,1,0,-1,0,-1,2,-2,1,0,1,1,-1,0,-2,-1,0,0,0,0,0,2,2,-1,-1,-1,-1,-1,1,1,-1,0,0,-1,0,0,1,-1,2,-1,-1,0,1,0,0,-1,-1,-1,-1};
			781: counter1_out = '{-2,0,0,0,1,1,0,-1,1,1,1,0,-1,-2,0,1,1,-1,0,0,1,1,1,-2,-1,0,0,1,0,0,-1,0,1,0,1,-1,-1,-1,0,0,2,1,0,-1,2,0,1,1,0,0,-1,0,1,0,-3,-1,0,1,-2,0,-1,-1,2,0,1,1,1,1,0,-2,1,0,1,0,-1,2,0,-1,-2,0,2,-1,2,1,-1,0,0,2,1,1,0,1,2,0,0,1,1,-1,-1,0};
			782: counter1_out = '{0,-1,1,0,0,1,-1,1,0,-2,0,1,-2,-1,-1,0,-1,1,0,0,-1,0,-2,-1,0,2,0,0,-1,0,0,0,0,-1,-2,0,-1,0,-1,0,0,-1,0,-1,2,1,0,1,1,-1,2,-1,1,1,1,0,0,1,0,-1,-1,0,-2,1,-2,0,0,1,0,0,1,1,0,-1,-1,-1,2,0,0,1,2,-1,0,0,-1,1,0,0,1,-1,0,1,1,1,1,0,-1,0,0,1};
			783: counter1_out = '{1,-1,1,1,-1,1,-1,-1,0,-1,-1,-1,1,-1,0,1,0,1,-1,-2,-1,0,-1,1,0,-1,-2,0,1,-2,-1,2,0,1,1,1,0,-1,0,1,-1,-1,1,0,-2,-1,1,0,1,0,-1,0,0,2,2,1,-2,0,0,0,1,-1,0,-1,2,1,0,1,2,0,1,2,0,0,1,0,0,1,0,1,0,0,-2,0,2,0,-1,-1,1,0,-1,0,0,-1,0,0,1,-1,-2,0};
			
		endcase
	end
	
	always_comb 
	// Combinational Block for counter2 matrix
	begin
		case (counter2)
			default: counter2_out = '{0,0,0,0,0,0,0,0,0,0};
			0: counter2_out = '{3,-2,-7,0,0,-2,-2,-5,2,7};
			1: counter2_out = '{2,-4,-4,1,-5,5,2,-1,6,-1};
			2: counter2_out = '{-2,-1,2,0,-4,-2,3,-3,-1,5};
			3: counter2_out = '{-3,1,7,1,-1,-1,1,0,-2,-5};
			4: counter2_out = '{-1,-2,-3,-1,-1,-4,1,0,-3,1};
			5: counter2_out = '{2,-1,1,-3,-6,-1,-2,1,2,4};
			6: counter2_out = '{2,-4,5,-2,-4,2,-1,-4,-2,4};
			7: counter2_out = '{1,3,1,0,0,-1,1,3,-3,-4};
			8: counter2_out = '{-1,0,1,5,1,4,-3,-4,-3,-4};
			9: counter2_out = '{-4,-2,2,-3,0,3,-4,2,0,0};
			10: counter2_out = '{0,-5,4,5,5,-3,-3,-2,0,-3};
			11: counter2_out = '{3,1,3,-3,-1,3,2,0,-7,-6};
			12: counter2_out = '{2,0,2,-3,0,2,-1,0,-3,1};
			13: counter2_out = '{-2,2,2,2,-4,-3,2,-2,1,3};
			14: counter2_out = '{-4,-4,3,2,-2,0,-2,-1,-2,-3};
			15: counter2_out = '{0,1,0,5,-2,-4,-1,2,-2,-4};
			16: counter2_out = '{-3,-2,3,-2,-1,2,-3,-3,2,1};
			17: counter2_out = '{-1,-2,-4,-2,6,4,-2,1,-4,-6};
			18: counter2_out = '{-1,-2,2,-6,-4,0,-1,-1,4,-1};
			19: counter2_out = '{2,0,-2,0,1,-2,-1,-3,5,0};
			20: counter2_out = '{-2,4,-9,-2,3,2,-1,5,-1,0};
			21: counter2_out = '{2,-5,-1,-2,2,0,-4,6,1,3};
			22: counter2_out = '{-1,0,2,5,-4,-4,-5,2,-5,-5};
			23: counter2_out = '{-1,2,2,-6,2,-2,0,5,3,-4};
			24: counter2_out = '{-1,2,-5,5,2,-1,-1,0,-4,-3};
			25: counter2_out = '{1,0,-2,-6,-3,2,0,2,4,-3};
			26: counter2_out = '{-3,-1,-5,1,-2,7,1,-2,-1,0};
			27: counter2_out = '{2,4,-1,0,6,-3,-1,-3,2,-3};
			28: counter2_out = '{-4,-3,-2,1,4,3,-6,-2,-9,4};
			29: counter2_out = '{3,2,3,-6,1,-4,-3,1,-1,-3};
			30: counter2_out = '{0,0,5,1,0,1,-2,0,2,-5};
			31: counter2_out = '{-4,0,-1,-3,2,3,-1,2,0,-2};
			32: counter2_out = '{-4,-2,3,-2,-2,3,0,-5,-2,3};
			33: counter2_out = '{-1,-2,-2,-2,-4,-1,-3,-2,2,0};
			34: counter2_out = '{-3,1,-1,3,0,-3,1,4,0,-3};
			35: counter2_out = '{3,5,-2,2,-2,0,1,-5,-2,1};
			36: counter2_out = '{-1,1,2,2,-2,-5,2,-3,-5,2};
			37: counter2_out = '{-5,0,-3,-5,-3,6,3,1,-8,-2};
			38: counter2_out = '{1,-2,1,6,0,-6,2,2,-2,-4};
			39: counter2_out = '{-5,0,-2,0,2,1,-1,-5,2,2};
			40: counter2_out = '{-3,2,-4,2,2,3,-1,1,-6,0};
			41: counter2_out = '{-3,-3,-4,2,4,2,-1,-4,4,-3};
			42: counter2_out = '{5,4,-1,-2,-3,1,2,-6,1,-4};
			43: counter2_out = '{-5,2,2,-4,-1,-1,3,2,-3,0};
			44: counter2_out = '{-6,-1,2,-4,-1,-2,1,-2,-2,3};
			45: counter2_out = '{-2,1,2,-2,-5,0,-3,0,0,4};
			46: counter2_out = '{1,2,1,-3,0,-1,3,2,-4,-3};
			47: counter2_out = '{-2,2,-3,-2,-4,6,5,3,-1,0};
			48: counter2_out = '{-1,-3,-2,7,1,-6,-2,-2,-2,-4};
			49: counter2_out = '{-4,0,4,1,-1,4,-8,-2,-5,-1};
			50: counter2_out = '{-1,1,-6,3,-1,-3,-2,3,-2,0};
			51: counter2_out = '{3,-1,-7,-5,0,-2,-6,4,-3,1};
			52: counter2_out = '{-3,1,3,-3,2,0,-3,2,0,0};
			53: counter2_out = '{0,1,0,-2,3,-1,1,3,-4,1};
			54: counter2_out = '{0,3,4,1,-1,6,-4,-3,-4,3};
			55: counter2_out = '{0,4,3,1,4,4,-2,-3,-5,-4};
			56: counter2_out = '{0,-1,-3,0,0,-3,0,1,4,-1};
			57: counter2_out = '{-2,-2,-3,-2,-2,5,4,2,-5,-1};
			58: counter2_out = '{2,3,-2,-2,4,2,-6,3,-1,0};
			59: counter2_out = '{-2,-2,2,-1,2,-2,-2,0,0,3};
			60: counter2_out = '{1,-3,0,2,-1,-1,1,0,-5,1};
			61: counter2_out = '{1,-2,-4,0,4,1,1,2,2,-4};
			62: counter2_out = '{-1,7,4,6,-5,-6,-1,0,-4,2};
			63: counter2_out = '{2,4,2,2,3,0,-3,-2,-1,-3};
			64: counter2_out = '{-4,-1,1,-3,-2,2,-1,3,1,-3};
			65: counter2_out = '{2,-1,3,-1,2,-1,0,-5,-7,5};
			66: counter2_out = '{-2,-2,-3,-6,-1,6,3,-1,1,0};
			67: counter2_out = '{-2,3,-3,-2,-1,4,1,6,-4,-1};
			68: counter2_out = '{1,-4,-2,5,1,-6,2,2,2,-3};
			69: counter2_out = '{1,0,-2,4,-2,4,-2,-3,-2,2};
			70: counter2_out = '{2,4,-2,-2,1,0,1,-6,0,-3};
			71: counter2_out = '{0,3,-2,1,2,0,1,0,-4,-1};
			72: counter2_out = '{-1,4,0,-2,7,-1,-3,1,-3,-6};
			73: counter2_out = '{1,0,-2,-4,0,-7,1,5,-1,-3};
			74: counter2_out = '{1,-1,2,3,-2,-3,3,-3,-5,-4};
			75: counter2_out = '{-3,-2,-5,4,-1,1,1,1,2,2};
			76: counter2_out = '{-5,1,-5,3,0,1,-6,-2,3,-1};
			77: counter2_out = '{0,0,-1,-6,-2,-4,-3,3,1,-1};
			78: counter2_out = '{3,1,-3,0,-3,2,-1,-3,-2,1};
			79: counter2_out = '{3,1,-3,3,0,-3,0,0,-2,-2};
			80: counter2_out = '{1,-2,6,-2,-2,-1,-1,-4,-2,3};
			81: counter2_out = '{2,1,0,0,-3,-1,-2,-2,1,4};
			82: counter2_out = '{4,2,1,1,-4,1,-3,2,0,-4};
			83: counter2_out = '{-1,-2,1,-2,-1,-1,1,0,2,2};
			84: counter2_out = '{-6,1,2,-2,-2,2,1,-1,-2,2};
			85: counter2_out = '{-5,-1,-5,-4,1,-5,-1,3,-3,1};
			86: counter2_out = '{0,-1,-1,3,-3,3,-2,4,-4,-6};
			87: counter2_out = '{-2,2,-5,-2,1,0,7,1,-3,-2};
			88: counter2_out = '{-3,-3,2,-3,-1,-3,4,2,3,-2};
			89: counter2_out = '{-4,2,-4,-3,-2,-1,5,-2,-2,4};
			90: counter2_out = '{-2,0,0,0,-7,2,3,0,2,-5};
			91: counter2_out = '{0,-1,-5,4,3,-2,0,3,0,0};
			92: counter2_out = '{0,-5,3,-3,-2,2,0,-1,0,3};
			93: counter2_out = '{2,-1,3,-2,4,-3,2,-3,-4,-4};
			94: counter2_out = '{-3,-3,-3,-1,-3,-1,-1,6,-2,-6};
			95: counter2_out = '{2,4,-3,2,2,-6,1,1,2,-2};
			96: counter2_out = '{-2,-1,4,2,-2,-4,-5,0,0,1};
			97: counter2_out = '{1,0,0,-4,5,0,1,-3,-3,-1};
			98: counter2_out = '{0,-3,-4,5,3,1,-1,-2,-3,4};
			99: counter2_out = '{1,-5,0,-3,-7,4,2,3,2,7};
		endcase
	end
	
endmodule 