module testbench();

timeunit 10ns;
timeprecision 1ns;

logic pixel, clk, reset, load, complete;
shortint result[0:9];

toplevel top0(.*);

always begin: CLOCK_GENERATION
	#1 clk = ~clk;
end

initial begin: CLOCK_INITIALIZATION
	clk = 0;
end



initial begin: TEST
#2 reset = 1;
load = 0;
#2 reset = 0;
load = 1;
#2 pixel = 0;
load = 0;

#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;

#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;

#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;

#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;

#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;

#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;

#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 1;
#2 pixel = 1;
#2 pixel = 1;
#2 pixel = 1;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;

#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 1;
#2 pixel = 1;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 1;
#2 pixel = 1;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;

#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 1;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 1;
#2 pixel = 1;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;

#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 1;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;

#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 1;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;

#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 1;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;

#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 1;
#2 pixel = 1;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;

#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 1;
#2 pixel = 1;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;

#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 1;
#2 pixel = 1;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;

#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 1;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;

#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 1;
#2 pixel = 1;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;

#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 1;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;

#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 1;
#2 pixel = 1;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;

#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 1;
#2 pixel = 1;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 1;
#2 pixel = 1;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;

#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 1;
#2 pixel = 1;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 1;
#2 pixel = 1;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;

#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 1;
#2 pixel = 1;
#2 pixel = 1;
#2 pixel = 1;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;

#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 1;
#2 pixel = 1;
#2 pixel = 1;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;

#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 1;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;

#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 1;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;

#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;

#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;

#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;
#2 pixel = 0;



end

endmodule
