// Top-level model

// Performs multiplication according to a state machine

module toplevel(input logic clk, reset, load, pixel, 
					output logic complete,
					output shortint result[0:9]);

	
	
	
	
	multiply_add multadd(.*);
	

	
endmodule