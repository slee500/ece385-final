// This is tthe top level file used in our final project

module final(input clk, );


LCD LCD0();


endmodule 