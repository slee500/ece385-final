
module nois (
	clk_clk,
	reset_reset_n,
	clk_27_clk);	

	input		clk_clk;
	input		reset_reset_n;
	output		clk_27_clk;
endmodule
